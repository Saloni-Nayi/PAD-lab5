�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   Ageq0X   Sexq1X   ChestPainTypeq2X	   RestingBPq3X   Cholesterolq4X	   FastingBSq5X
   RestingECGq6X   MaxHRq7X   ExerciseAnginaq8X   Oldpeakq9X   ST_Slopeq:etq;bX   n_features_in_q<KX
   n_outputs_q=KX   classes_q>h"h#K �q?h%�q@RqA(KK�qBh)X   i8qC���qDRqE(KX   <qFNNNJ����J����K tqGb�C               qHtqIbX
   n_classes_qJKX   base_estimator_qKhX   estimators_qL]qM(h)�qN}qO(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h<Kh=Kh>h"h#K �qPh%�qQRqR(KK�qSh)X   f8qT���qURqV(KhFNNNJ����J����K tqWb�C              �?qXtqYbhJcnumpy.core.multiarray
scalar
qZhEC       q[�q\Rq]X   max_features_q^KX   tree_q_csklearn.tree._tree
Tree
q`Kh"h#K �qah%�qbRqc(KK�qdhE�C       qetqfbK�qgRqh}qi(hKX
   node_countqjMSX   nodesqkh"h#K �qlh%�qmRqn(KMS�qoh)X   V56qp���qqRqr(Kh-N(X
   left_childqsX   right_childqtX   featurequX	   thresholdqvX   impurityqwX   n_node_samplesqxX   weighted_n_node_samplesqytqz}q{(hsh)X   i8q|���q}Rq~(KhFNNNJ����J����K tqbK �q�hth~K�q�huh~K�q�hvhVK�q�hwhVK �q�hxh~K(�q�hyhVK0�q�uK8KKtq�b�B(J         �                    �?j8je3�?�           ��@       #                    �?�}�	���?           �y@                           @I@^n����?'             N@       	                     E@�q�q�?             2@                           �B@����X�?             @                           W@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @
                           �H@�C��2(�?
             &@������������������������       �                      @                          @N@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?       "                    �P@r�q��?             E@                           U@�p ��?            �D@                           @M@      �?             @@                           �L@�KM�]�?             3@                           @J@��S�ۿ?	             .@                           C@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@                           P@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@       !                    @O@X�<ݚ�?             "@                           �U@�q�q�?             @                          `U@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?$       o                   @O@�g���E�?�             v@%       l                    �R@�BѶ�n�?�            �m@&       )                    @3e��?�            `m@'       (                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @*       O                   �I@��ϭ�*�?�             m@+       <                    �I@�}�+r��?l            `e@,       3                   �B@�KM�]�?             C@-       0                     I@z�G�z�?	             .@.       /                    �D@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@1       2                   �?@�q�q�?             @������������������������       �                     �?������������������������       �                      @4       ;                   @G@�nkK�?             7@5       6                   �F@��S�ۿ?             .@������������������������       �                     @7       :                     H@ףp=
�?             $@8       9                    @F@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @=       N                   @B@0�!F��?W            �`@>       K                   �A@ ��Ou��?1            �S@?       @                    @L@hA� �?,            �Q@������������������������       �                     :@A       D                    �L@t��ճC�?             F@B       C                    5@      �?             @������������������������       �                     @������������������������       �                     �?E       J                    .@P���Q�?             D@F       G                    +@"pc�
�?             &@������������������������       �                     @H       I                    �N@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     =@L       M                    @L@      �?              @������������������������       �      �?             @������������������������       �                     @������������������������       �        &            �K@P       S                   @J@L=�m��?%            �N@Q       R                     L@�q�q�?             (@������������������������       �                      @������������������������       �                     @T       a                   �L@؇���X�?            �H@U       `                   @L@�>4և��?             <@V       W                   �J@PN��T'�?             ;@������������������������       �                      @X       [                   @K@�J�4�?             9@Y       Z                    �O@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @\       ]                    �F@؇���X�?	             ,@������������������������       �                     @^       _                     M@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?b       c                   @M@�����?             5@������������������������       �                     @d       k                    �M@؇���X�?             ,@e       f                   @N@$�q-�?             *@������������������������       �                     @g       j                    �I@r�q��?             @h       i                    �G@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?m       n                    B@      �?              @������������������������       �                     �?������������������������       �                     �?p       �                    Y@r�����?E            �\@q       �                   �P@">�֕�?A            @Z@r       �                   �P@�eP*L��?            �@@s       x                    �H@     ��?             @@t       w                    @F@z�G�z�?             $@u       v                     D@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @y       z                    @I@���!pc�?             6@������������������������       �                     @{       |                    @J@�����?             3@������������������������       �                      @}       �                   @P@������?             1@~                            P@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �K@d}h���?	             ,@������������������������       �                      @�       �                    �L@      �?             (@������������������������       �                     �?�       �                    @M@"pc�
�?             &@������������������������       �                     @�       �                    �M@      �?              @������������������������       �                     �?�       �                     P@؇���X�?             @������������������������       �                     @�       �                    `P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �M@      �?,             R@�       �                   `R@��X��?%             L@�       �                   `Q@d}h���?             ,@�       �                    @I@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �D@X�Cc�?             E@�       �                    �B@@4և���?
             ,@�       �                    �A@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                   �R@      �?             <@������������������������       �                     @�       �                    �F@� �	��?             9@������������������������       �                     @�       �                    @J@�q�q�?             5@������������������������       �                     "@�       �                   �U@�q�q�?             (@�       �                   �R@�<ݚ�?             "@������������������������       �                     �?�       �                   �S@      �?              @�       �                    @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     0@�       �                    �D@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                   @I@"\�����?�             t@�       �                    @K@�q�q�?,            @Q@�       �                    �H@������?             1@�       �                    �?���|���?	             &@������������������������       �                     @�       �                   �E@�q�q�?             @�       �                    7@�q�q�?             @������������������������       �                     �?�       �                    �G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?���B���?             J@�       �                    C@���Q��?             $@�       �                    �L@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                     P@�����?             E@�       �                    �?(;L]n�?             >@������������������������       �                     @�       �                    B@�nkK�?             7@�       �                    :@�����H�?             "@������������������������       �                     @�       �                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@�       �                    �?      �?             (@������������������������       �                     �?�       �                    �P@���!pc�?             &@������������������������       �                     �?�       �                    @z�G�z�?             $@�       �                    �Q@�<ݚ�?             "@������������������������       �                     @�       �                    @R@�q�q�?             @�       �                    A@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �?:]���?�            �o@�       �                   �W@���;QU�?/            @R@�       �                    �?@3����?$             K@������������������������       �                     A@�       �                    @I@P���Q�?             4@�       �                   `P@ףp=
�?             $@������������������������       �                     @�       �                     H@z�G�z�?             @������������������������       �                     @�       �                   �R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                    @G@���y4F�?             3@������������������������       �                     &@�       �                    @      �?              @�       �                    @I@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   �K@���Z�?u            �f@������������������������       �                      @�       B                   @�μ���?t            @f@�       1                  �W@��ɉ��?e            �c@�                          @K@��Xk�?I             \@�       �                    @B@�j��b�?)            �M@�       �                    R@���Q��?             @������������������������       �                     �?�       �                    �A@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    W@�>����?$             K@�       �                   `P@`'�J�?"            �I@�       �                    @H@      �?
             0@������������������������       �                      @�       �                    @I@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                    �A@                          �?�q�q�?             @������������������������       �                      @������������������������       �                     �?      "                   @M@Fmq��?             �J@                         @L@��
ц��?            �C@                        �M@      �?
             8@������������������������       �                      @                         �K@�X����?	             6@      	                  �P@ҳ�wY;�?             1@������������������������       �                     @
                         R@���Q��?             $@������������������������       �                     @                         �?�q�q�?             @������������������������       �                     @������������������������       �                      @                        �S@z�G�z�?             @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        `R@���Q��?	             .@                         �?      �?             @                         Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                         �?�eP*L��?             &@                        @T@�q�q�?             @������������������������       �                      @������������������������       �                     �?                         �L@      �?              @������������������������       �                     �?       !                   V@և���X�?             @������������������������       �                     �?������������������������       ��q�q�?             @#      *                   �O@d}h���?             ,@$      )                   @N@�����H�?	             "@%      &                  �P@z�G�z�?             @������������������������       �                      @'      (                   �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @+      ,                   �?���Q��?             @������������������������       �                      @-      .                   �P@�q�q�?             @������������������������       �                     �?/      0                  �R@      �?              @������������������������       �                     �?������������������������       �                     �?2      3                  �X@�����H�?            �F@������������������������       �        	             0@4      9                   �?д>��C�?             =@5      6                   �I@��S�ۿ?	             .@������������������������       �                     "@7      8                  �[@r�q��?             @������������������������       �                     @������������������������       �                     �?:      A                  �Z@����X�?
             ,@;      @                   �L@���Q��?             $@<      =                   Y@      �?              @������������������������       �                     @>      ?                   @G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @C      R                   �O@և���X�?             5@D      M                  �U@�q�q�?             2@E      J                   �N@"pc�
�?             &@F      I                  �P@�����H�?             "@G      H                   @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @K      L                  �N@      �?              @������������������������       �                     �?������������������������       �                     �?N      Q                  @Z@և���X�?             @O      P                   �L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KMSKK�q�hV�B0       Ps@     �z@      U@     �t@      3@     �D@      (@      @       @      @       @       @               @       @                      @      $@      �?       @               @      �?      �?      �?      �?              @     �A@      @     �A@       @      >@       @      1@      �?      ,@      �?      @      �?                      @              "@      �?      @      �?                      @              *@      @      @      @       @      �?       @      �?                       @      @                      @      �?             @P@     �q@      7@     �j@      6@     �j@       @      �?              �?       @              4@     �j@      "@     @d@      @      A@      @      (@      �?      &@      �?                      &@       @      �?              �?       @              �?      6@      �?      ,@              @      �?      "@      �?      @              @      �?                      @               @      @      `@      @     @R@      @     �P@              :@      @     �D@      �?      @              @      �?               @      C@       @      "@              @       @       @               @       @                      =@       @      @       @       @              @             �K@      &@      I@      @       @               @      @              @      E@      @      7@      @      7@               @      @      5@       @      "@              "@       @               @      (@              @       @      @       @                      @      �?               @      3@              @       @      (@      �?      (@              @      �?      @      �?       @               @      �?                      @      �?              �?      �?              �?      �?              E@     @R@     �@@      R@      .@      2@      ,@      2@       @       @      @       @      @                       @      @              @      0@              @      @      *@       @              @      *@      �?       @               @      �?              @      &@               @      @      "@      �?               @      "@              @       @      @      �?              �?      @              @      �?       @      �?                       @      �?              2@      K@      2@      C@      @      &@      @      @      @                      @              @      .@      ;@      �?      *@      �?      @              @      �?                      "@      ,@      ,@      @              &@      ,@      @              @      ,@              "@      @      @      @       @              �?      @      �?       @      �?              �?       @              @                      @              0@      "@      �?              �?      "@              l@     @X@      7@      G@      *@      @      @      @      @               @      @       @      �?      �?              �?      �?      �?                      �?              @      @              $@      E@      @      @       @      @       @                      @      @              @      C@      �?      =@              @      �?      6@      �?       @              @      �?      @      �?                      @              ,@      @      "@              �?      @       @      �?               @       @       @      @              @       @      @       @      �?              �?       @                      @              �?     @i@     �I@      Q@      @     �J@      �?      A@              3@      �?      "@      �?      @              @      �?      @              �?      �?              �?      �?              $@              .@      @      &@              @      @      @      @              @      @              �?             �`@      G@               @     �`@      F@     @_@      @@     @U@      ;@     �J@      @      @       @              �?      @      �?      @                      �?      I@      @     �H@       @      ,@       @       @              @       @               @      @             �A@              �?       @               @      �?              @@      5@      5@      2@      .@      "@               @      .@      @      &@      @      @              @      @              @      @       @      @                       @      @      �?      �?      �?      �?                      �?      @              @      "@      �?      @      �?       @      �?                       @              �?      @      @       @      �?       @                      �?      @      @              �?      @      @      �?               @      @      &@      @       @      �?      @      �?       @               @      �?       @                      �?      @              @       @       @              �?       @              �?      �?      �?              �?      �?              D@      @      0@              8@      @      ,@      �?      "@              @      �?      @                      �?      $@      @      @      @      @       @      @              �?       @      �?                       @               @      @              "@      (@      @      (@       @      "@      �?       @      �?       @      �?                       @              @      �?      �?              �?      �?              @      @      @      �?      @                      �?               @      @        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hKhjM_hkh"h#K �q�h%�q�Rq�(KM_�q�hr�B�L         �                   �M@4�5����?�           ��@       %                    �?�������?�            �s@                           �M@^H���+�?            �B@                           �J@� �	��?             9@                          �H@������?             .@                           �?�����H�?             "@                          �:@z�G�z�?             @������������������������       �                     �?	       
                    �G@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     @                          @K@      �?             @������������������������       �                      @                           �?      �?             @                            F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                            L@�z�G��?             $@������������������������       �                     @                            @���Q��?             @                           �L@      �?             @������������������������       �                     �?                          @G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                           �N@r�q��?	             (@������������������������       �                     @                            �?�<ݚ�?             "@������������������������       �                     �?!       "                    �Q@      �?              @������������������������       �                     @#       $                    `R@�q�q�?             @������������������������       �                     �?������������������������       �                      @&                           �?r ��*�?�            �q@'       |                    �R@�KM�]�?�             j@(       {                     P@�θV�?�            �i@)       *                    @�y��*�?n            �e@������������������������       �                     �?+       <                   @@@��㨇,�?m            �e@,       -                    +@      �?#             P@������������������������       �                     ,@.       1                    .@HP�s��?             I@/       0                    �N@      �?             @������������������������       �                      @������������������������       �                      @2       3                   �:@�nkK�?             G@������������������������       �                     5@4       9                    �O@HP�s��?             9@5       6                    �L@�nkK�?             7@������������������������       �                     ,@7       8                    =@�����H�?             "@������������������������       �      �?              @������������������������       �                     @:       ;                   �=@      �?              @������������������������       �                     �?������������������������       �                     �?=       ^                    @L@>����?J            @[@>       Q                    �I@�θV�?/            @Q@?       @                   @A@6YE�t�?            �@@������������������������       �                     �?A       D                    �F@      �?             @@B       C                   �D@��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@E       P                   �K@@�0�!��?             1@F       O                    �G@      �?             0@G       L                    @G@z�G�z�?             $@H       I                   @E@r�q��?             @������������������������       �                     @J       K                   @H@�q�q�?             @������������������������       �                     �?������������������������       �                      @M       N                   @I@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?R       S                    @J@�X�<ݺ?             B@������������������������       �                     @T       W                    �J@ 	��p�?             =@U       V                    D@؇���X�?             @������������������������       �                     �?������������������������       �                     @X       Y                    @K@���7�?             6@������������������������       �                      @Z       ]                    �K@@4և���?
             ,@[       \                   @B@�����H�?             "@������������������������       �      �?              @������������������������       �                     @������������������������       �                     @_       z                   �L@R���Q�?             D@`       k                    �M@���"͏�?            �B@a       b                   @B@��Q��?             4@������������������������       �                     @c       d                   @I@������?             1@������������������������       �                     "@e       j                    @M@      �?              @f       i                    �L@�q�q�?             @g       h                   @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @l       q                    @N@�t����?             1@m       n                    D@z�G�z�?             @������������������������       �                     @o       p                    I@      �?              @������������������������       �                     �?������������������������       �                     �?r       s                   �E@�8��8��?	             (@������������������������       �                     @t       u                    @O@z�G�z�?             @������������������������       �                     �?v       y                    �O@      �?             @w       x                   @G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                    �@@}       ~                    B@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @K@X~�pX��?1            @R@�       �                    �J@�q�q�?             2@�       �                     F@�eP*L��?	             &@������������������������       �                      @�       �                   @E@�q�q�?             "@������������������������       �                     @�       �                   �F@      �?             @������������������������       �                      @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?%            �K@�       �                    @L@�z�G��?             $@������������������������       �                     �?�       �                   �K@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    @:	��ʵ�?            �F@�       �                   �E@��G���?            �B@�       �                    @R@�	j*D�?
             *@�       �                     N@�����H�?             "@�       �                    @M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �?@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    J@      �?             8@�       �                    �M@�X�<ݺ?             2@�       �                    @M@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@�       �                   �K@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    K@      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?l�?���?�            �y@�       �                    �?"pc�
�?B            @^@�       �                   �T@��+��?            �B@�       �                    Q@���y4F�?             3@�       �                     M@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �S@�r����?	             .@������������������������       �                      @�       �                    �O@����X�?             @������������������������       �                     @������������������������       �                      @�       �                   �V@�<ݚ�?             2@�       �                   �U@      �?             0@�       �                    U@      �?              @������������������������       �                     @�       �                    �L@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    �?h�����?0             U@������������������������       �                    �D@�       �                    @Du9iH��?            �E@�       �                   �T@ >�֕�?            �A@�       �                     I@�<ݚ�?             "@�       �                    S@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     :@�       �                   @R@      �?              @�       �                    Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       *                   @L@D�]�+��?�            `r@�                          @J@��/���?�            `j@�       �                    �? �D^��?d            @d@�       �                   �R@�y(dD�?%            @P@�       �                   @N@����X�?             5@������������������������       �                     @�       �                    @D@r�q��?             2@������������������������       �                     �?�       �                   `P@�t����?
             1@������������������������       �                     @�       �                   �P@r�q��?             (@�       �                     H@      �?              @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @�       �                   @[@"pc�
�?             F@�       �                   �U@$�q-�?            �C@������������������������       �        	             1@�       �                    V@��2(&�?             6@�       �                    �G@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �W@ףp=
�?             4@������������������������       �                     "@�       �                    �D@"pc�
�?             &@������������������������       �                     @�       �                   `X@�q�q�?             @�       �                    @G@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @�                          @L� P?)�??            @X@�       �                    �?J� ��w�?<             W@�       �                   �W@8�Z$���?              J@�       �                    W@l��
I��?             ;@�       �                     G@      �?             8@�       �                    �@@ҳ�wY;�?             1@������������������������       �                     @�       �                    �B@և���X�?
             ,@������������������������       �                     @�       �                    �E@���!pc�?             &@������������������������       �                     @�       �                    Q@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     9@                          �F@z�G�z�?             D@������������������������       �                     8@                        �R@     ��?             0@������������������������       �                      @                        �Y@X�Cc�?
             ,@                        �S@      �?	             (@                         @G@      �?             @������������������������       �                      @������������������������       �                      @	      
                  �X@      �?              @������������������������       �                     @                         @H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                         @F@z�G�z�?             @                         �C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @      )                  @[@���c�H�?            �H@      (                   �K@�㙢�c�?             G@      '                  `T@� ��1�?            �D@                         �J@r֛w���?             ?@                        �P@���!pc�?             &@                         �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                         P@      �?             4@������������������������       �                     "@                         �P@�eP*L��?             &@������������������������       �                     �?!      &                   �?���Q��?             $@"      %                   �?؇���X�?             @#      $                  �R@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@������������������������       �                     @������������������������       �                     @+      @                   �?NP�<��?4            �T@,      9                  �P@      �?             D@-      0                  @P@������?             .@.      /                   �O@      �?              @������������������������       �                     �?������������������������       �                     �?1      4                   �M@�θ�?	             *@2      3                   @M@      �?             @������������������������       �                      @������������������������       �                      @5      6                    P@�����H�?             "@������������������������       �                     @7      8                   `P@�q�q�?             @������������������������       �                     �?������������������������       �                      @:      ?                  �R@`2U0*��?             9@;      >                   �M@      �?              @<      =                   R@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        
             1@A      ^                  �U@X��ʑ��?            �E@B      ]                  `U@h+�v:�?             A@C      N                   �M@П[;U��?             =@D      G                   �L@���!pc�?             &@E      F                  �P@z�G�z�?             @������������������������       �                     �?������������������������       �                     @H      I                   �?�q�q�?             @������������������������       �                     �?J      M                   @M@z�G�z�?             @K      L                  @R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @O      \                   `Q@�E��ӭ�?             2@P      [                    Q@     ��?
             0@Q      Z                  �T@������?	             .@R      S                  �P@8�Z$���?             *@������������������������       �                     @T      U                  `Q@����X�?             @������������������������       �                     �?V      W                   @r�q��?             @������������������������       �                     �?X      Y                   @O@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@q�tq�bh�h"h#K �q�h%�q�Rq�(KM_KK�q�hV�B�       �t@     y@     @Q@     @o@      8@      *@      ,@      &@      &@      @       @      �?      @      �?      �?              @      �?      �?               @      �?      @              @      @               @      @      �?       @      �?              �?       @              �?              @      @              @      @       @       @       @              �?       @      �?              �?       @              �?              $@       @      @              @       @              �?      @      �?      @               @      �?              �?       @             �F@     �m@      6@     `g@      5@     @g@      5@      c@      �?              4@      c@      @      N@              ,@      @      G@       @       @               @       @               @      F@              5@       @      7@      �?      6@              ,@      �?       @      �?      �?              @      �?      �?              �?      �?              0@     @W@      @      O@      @      <@      �?              @      <@      �?      ,@      �?                      ,@      @      ,@       @      ,@       @       @      �?      @              @      �?       @      �?                       @      �?      @              @      �?                      @      �?               @      A@              @       @      ;@      �?      @      �?                      @      �?      5@               @      �?      *@      �?       @      �?      �?              @              @      "@      ?@      "@      <@      @      *@      @              @      *@              "@      @      @       @      @       @      �?       @                      �?              @       @               @      .@      �?      @              @      �?      �?      �?                      �?      �?      &@              @      �?      @              �?      �?      @      �?       @      �?                       @              �?              @             �@@      �?      �?              �?      �?              7@      I@      (@      @      @      @       @              @      @              @      @      @       @              �?      @              @      �?              @              &@      F@      @      @      �?               @      @              @       @               @     �B@      @      >@      @      "@      �?       @      �?      �?              �?      �?                      @      @      �?              �?      @              @      5@      �?      1@      �?      @              @      �?                      &@       @      @       @                      @      �?      @              @      �?             �p@     �b@     �X@      6@      2@      3@      @      .@       @       @       @                       @       @      *@               @       @      @              @       @              ,@      @      ,@       @      @       @      @              @       @      @                       @       @                       @     @T@      @     �D@              D@      @     �@@       @      @       @      @       @      @                       @      @              :@              @      �?      �?      �?      �?                      �?      @             �d@      `@     `a@      R@     @Y@     �N@      7@      E@      .@      @              @      .@      @              �?      .@       @      @              $@       @      @       @      @              �?       @      @               @      B@      @      B@              1@      @      3@      �?      �?      �?                      �?       @      2@              "@       @      "@              @       @      @       @       @       @                       @               @      @             �S@      3@     @S@      .@      F@       @      3@       @      2@      @      &@      @      @               @      @              @       @      @      @               @      @       @                      @      @              �?       @      �?                       @      9@             �@@      @      8@              "@      @               @      "@      @      "@      @       @       @       @                       @      @      �?      @               @      �?       @                      �?               @      �?      @      �?      �?              �?      �?                      @      C@      &@      C@       @     �@@       @      7@       @       @      @       @      @              @       @              @              .@      @      "@              @      @              �?      @      @      @      �?       @      �?              �?       @              @                      @      $@              @                      @      :@     �L@      @     �A@      @      &@      �?      �?              �?      �?              @      $@       @       @               @       @              �?       @              @      �?       @      �?                       @      �?      8@      �?      @      �?      @              @      �?                      @              1@      5@      6@      5@      *@      0@      *@      @       @      �?      @      �?                      @       @      @      �?              �?      @      �?      �?              �?      �?                      @      *@      @      &@      @      &@      @      &@       @      @              @       @              �?      @      �?      �?              @      �?              �?      @                       @              �?       @              @                      "@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hKhjM}hkh"h#K �q�h%�q�Rq�(KM}�q�hr�BXS         �                   �M@p�Vv���?�           ��@                           �?�dG��?�            �t@                           �M@v�X��?             F@                           @J@*;L]n�?             >@                           J@�GN�z�?             6@                           �G@�t����?             1@������������������������       �                     @                          �A@"pc�
�?             &@	       
                    �H@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @                           �H@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     ,@       '                    �I@�k�'7��?�            �q@                           �?     8�?(             P@                           �F@��Y��]�?            �D@������������������������       �        
             4@                           @G@���N8�?             5@                          @E@؇���X�?             @������������������������       �                     @                          @H@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@       &                    �H@�LQ�1	�?             7@       %                    @z�G�z�?
             .@                            �?؇���X�?	             ,@������������������������       �                     @!       "                    7@      �?              @������������������������       �                      @#       $                    @G@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @(       m                    �?�K��E/�?�            �k@)       l                     P@ w���?v            �d@*       A                   �;@ȖLy�r�?b            �`@+       <                    :@z�G�z�?            �A@,       -                    +@ȵHPS!�?             :@������������������������       �                     $@.       ;                   �7@     ��?             0@/       6                    5@���!pc�?
             &@0       5                    .@؇���X�?             @1       2                    �N@�q�q�?             @������������������������       �                     �?3       4                    @O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @7       8                    @K@      �?             @������������������������       �                     �?9       :                    @N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @=       >                    @L@X�<ݚ�?             "@������������������������       �                      @?       @                    �L@և���X�?             @������������������������       �                      @������������������������       ����Q��?             @B       [                    @O@�"P��?I            �X@C       R                   �I@xdQ�m��?;            @T@D       I                    �J@��ɉ�?-            @P@E       H                    E@ףp=
�?             $@F       G                   �A@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @J       K                    �L@ �Jj�G�?&            �K@������������������������       �                     8@L       Q                   @B@�g�y��?             ?@M       P                    �M@�8��8��?	             (@N       O                   �@@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                     3@S       T                    @L@     ��?             0@������������������������       �                     @U       V                   �J@�z�G��?             $@������������������������       �                      @W       X                   @L@      �?              @������������������������       �                     @Y       Z                    @M@      �?             @������������������������       �                     @������������������������       �                     �?\       c                    F@r�q��?             2@]       ^                    �O@�C��2(�?             &@������������������������       �                     @_       `                   �=@r�q��?             @������������������������       �                     @a       b                   �A@�q�q�?             @������������������������       �                     �?������������������������       �                      @d       e                   @G@����X�?             @������������������������       �                     �?f       k                   �K@r�q��?             @g       h                    �O@�q�q�?             @������������������������       �                     �?i       j                   �I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                    �@@n       �                   �K@������?'             K@o       �                   @H@��[�p�?"            �G@p       �                   �C@��R[s�?            �A@q       v                   �0@R���Q�?             4@r       s                    �N@�q�q�?             @������������������������       �                     �?t       u                    $@      �?              @������������������������       �                     �?������������������������       �                     �?w       x                   �:@�t����?             1@������������������������       �                     @y       �                    @z�G�z�?	             $@z       }                    �?      �?              @{       |                     L@�q�q�?             @������������������������       �                     �?������������������������       �                      @~                           �N@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @���Q��?	             .@�       �                    �P@      �?             (@�       �                    �?      �?              @������������������������       �                     �?�       �                     L@����X�?             @������������������������       �                     �?�       �                    �M@r�q��?             @�       �                    @M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�8��8��?             (@������������������������       �                     @�       �                    @r�q��?             @�       �                    J@�q�q�?             @������������������������       �                     �?�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @K@և���X�?             @������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                     �?�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�                          �?���Q��?           Py@�       �       	             �?�`⯛��?c            �c@�       �                    `P@H�V�e��?             A@�       �                   �X@     ��?             @@�       �                   �S@��� ��?             ?@������������������������       �        	             .@�       �                    �O@      �?             0@�       �                    @M@z�G�z�?
             .@�       �                     F@�q�q�?             @������������������������       �                     @�       �                   �T@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �N@�����H�?             "@������������������������       �                     @�       �                    U@r�q��?             @�       �                   `T@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    P@ҐϿ<��?M            �^@�       �                   @O@�n_Y�K�?	             *@�       �                    �G@      �?             @������������������������       �                      @�       �                    �J@      �?             @�       �                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                     L@����X�?             @������������������������       �                     @�       �                     P@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �M@����x�?D            @[@�       �                    �D@t�����?4             U@�       �                    R@ףp=
�?             4@�       �                     D@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �B@�IєX�?
             1@�       �                    V@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                   �Q@     ��?(             P@�       �                     H@l��
I��?             ;@�       �                    Q@���Q��?             @�       �                    @F@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                     M@�GN�z�?             6@�       �                     L@�t����?             1@�       �                    @K@z�G�z�?             $@�       �                    �I@�����H�?             "@�       �                   `P@r�q��?             @������������������������       �                      @������������������������       �      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �P@���Q��?             @������������������������       �      �?             @������������������������       �                     �?�       �                   �U@��J�fj�?            �B@�       �                   �S@$��m��?             :@�       �                    �F@      �?             0@������������������������       �                      @�       �                    �I@և���X�?
             ,@������������������������       �                     @�       �                    �K@�eP*L��?             &@�       �                   �R@����X�?             @������������������������       �                     @�       �                    @K@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �R@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?�       �                    U@ףp=
�?             $@�       �                   `T@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   `[@���|���?	             &@�       �                    �E@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                      @�                         �P@H%u��?             9@�       �                     P@�q�q�?             "@������������������������       �                     @�                           `P@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@                         �?��-�?�             o@                         @H@�����?,            �P@������������������������       �                    �@@                         �I@l��\��?             A@                        @U@���Q��?             @                         �H@�q�q�?             @	      
                  �Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         R@XB���?             =@                         Q@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     3@      F                   @K@����X�?t            �f@      A                   @��G���?F            �[@                          �E@�`�=	�?@            �Y@                         Q@�nkK�?             G@                         �B@      �?             @������������������������       �                     �?������������������������       �                     @                         �?�Ń��̧?             E@                        �V@���7�?             6@                        �T@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@������������������������       �                     4@!      4                   @I@���y4F�?"            �L@"      3                   @H@b�h�d.�?            �A@#      $                  �Q@�θ�?             :@������������������������       �                     @%      0                   �G@�����?
             3@&      +                   �?      �?             0@'      *                   �F@�z�G��?             $@(      )                  �U@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @,      /                   @G@r�q��?             @-      .                   �F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @1      2                  �V@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@5      :                   �?���!pc�?             6@6      7                   �J@�8��8��?             (@������������������������       �                      @8      9                  @[@      �?             @������������������������       �                     @������������������������       �                     �?;      <                  �Q@      �?             $@������������������������       �                     @=      >                  @S@����X�?             @������������������������       �                     @?      @                   X@      �?             @������������������������       �                      @������������������������       �                      @B      E                  @Z@      �?              @C      D                  �Y@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @G      |                    Q@R_u^|�?.            �Q@H      q                   �N@j���� �?-             Q@I      d                   @M@~|z����?#            �J@J      c                   @���Q��?            �A@K      R                   �K@�4�����?             ?@L      O                   �?"pc�
�?             &@M      N                   R@؇���X�?             @������������������������       �                     �?������������������������       �                     @P      Q                  �Q@      �?             @������������������������       �                     @������������������������       �                     �?S      X                   �L@���Q��?             4@T      W                  `S@�q�q�?             "@U      V                  �P@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @Y      Z                   Q@�eP*L��?             &@������������������������       �                      @[      b                  �W@�q�q�?             "@\      ]                  �T@      �?              @������������������������       �                      @^      a                   V@�q�q�?             @_      `                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     @e      n                   @N@b�2�tk�?             2@f      g                   �?�	j*D�?	             *@������������������������       �                     @h      m                   @ףp=
�?             $@i      l                  @P@؇���X�?             @j      k                  @N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @o      p                   @���Q��?             @������������������������       �                     @������������������������       �                      @r      s                  @N@z�G�z�?
             .@������������������������       �                     �?t      {                  @W@؇���X�?	             ,@u      v                   �P@$�q-�?             *@������������������������       �                     "@w      z                   @      �?             @x      y                   S@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KM}KK�q�hV�B�       @t@     �y@     @T@      o@      ?@      *@      1@      *@      1@      @      .@       @      @              "@       @      @       @               @      @              @               @      @       @                      @               @      ,@              I@     `m@      5@     �E@      �?      D@              4@      �?      4@      �?      @              @      �?      @      �?                      @              ,@      4@      @      (@      @      (@       @      @              @       @       @              @       @      @                       @              �?       @              =@      h@      .@      c@      .@     �]@      @      <@      @      7@              $@      @      *@      @       @      �?      @      �?       @              �?      �?      �?      �?                      �?              @       @       @              �?       @      �?       @                      �?              @      @      @               @      @      @       @               @      @       @     �V@      @      S@       @     �O@      �?      "@      �?      @              @      �?                      @      �?      K@              8@      �?      >@      �?      &@      �?       @               @      �?                      "@              3@      @      *@              @      @      @       @              �?      @              @      �?      @              @      �?              @      .@      �?      $@              @      �?      @              @      �?       @      �?                       @       @      @      �?              �?      @      �?       @              �?      �?      �?              �?      �?                      @             �@@      ,@      D@      $@     �B@      "@      :@      @      1@      �?       @              �?      �?      �?              �?      �?               @      .@              @       @       @       @      @      �?       @      �?                       @      �?      @      �?                      @               @      @      "@      @      @       @      @              �?       @      @      �?              �?      @      �?       @               @      �?                      @      @                      @      �?      &@              @      �?      @      �?       @              �?      �?      �?      �?                      �?              @      @      @       @               @      @      �?              �?      @              @      �?             `n@     @d@     �H@     �Z@      @      ;@      @      ;@      @      ;@              .@      @      (@      @      (@       @      @              @       @      �?              �?       @              �?       @              @      �?      @      �?      �?              �?      �?                      @      �?              �?               @              E@      T@       @      @      @      @               @      @      �?      �?      �?      �?                      �?       @              @       @      @               @       @               @       @              A@     �R@      ?@     �J@       @      2@      �?       @               @      �?              �?      0@      �?      @              @      �?                      $@      =@     �A@       @      3@      @       @      @      �?              �?      @                      �?      @      1@       @      .@       @       @      �?       @      �?      @               @      �?      @              @      �?                      @      @       @      @      �?              �?      5@      0@      1@      "@       @       @       @              @       @              @      @      @      @       @      @               @       @               @       @              �?      @      �?       @              �?      "@      �?      @      �?      @                      �?      @              @      @       @      @       @                      @       @              @      6@      @      @              @      @      �?      @                      �?              0@     @h@     �K@      P@      @     �@@              ?@      @      @       @      �?       @      �?      �?      �?                      �?              �?       @              <@      �?      "@      �?      "@                      �?      3@             @`@      J@     �V@      5@     @V@      ,@      F@       @      @      �?              �?      @             �D@      �?      5@      �?      @      �?      @                      �?      ,@              4@             �F@      (@      =@      @      4@      @      @              *@      @      (@      @      @      @      @      @              @      @              @              @      �?       @      �?       @                      �?      @              �?       @      �?                       @      "@              0@      @      &@      �?       @              @      �?      @                      �?      @      @      @               @      @              @       @       @       @                       @      �?      @      �?      @              @      �?                      @      D@      ?@      D@      <@      <@      9@      5@      ,@      5@      $@      "@       @      @      �?              �?      @              @      �?      @                      �?      (@       @      @      @       @      @       @                      @      @              @      @               @      @      @      @       @       @              @       @       @      �?              �?       @               @      �?              �?              @      @      &@      @      "@      @              �?      "@      �?      @      �?      �?              �?      �?                      @              @      @       @      @                       @      (@      @              �?      (@       @      (@      �?      "@              @      �?       @      �?              �?       @              �?                      �?              @q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       qنq�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hKhjMYhkh"h#K �q�h%�q�Rq�(KMY�q�hr�BxK         D       	             �?U�ք�?�           ��@       '                    �?�Q����?i             d@       &                   �X@     ��?%             P@                           �J@������?#             N@                          �V@
;&����?             7@                          �M@և���X�?             5@                           �G@���|���?             &@������������������������       �                     @	       
                    �H@      �?              @������������������������       �                     @                          @F@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @                           �D@z�G�z�?             $@������������������������       �                     �?                           R@�����H�?             "@������������������������       �                     @                            I@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                          �N@������?            �B@                          @L@���!pc�?	             &@                          �E@z�G�z�?             $@������������������������       �                     @                           �P@����X�?             @                          �G@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?        !                    �N@ ��WV�?             :@������������������������       �                     *@"       #                    U@$�q-�?             *@������������������������       �                     @$       %                   �V@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @(       -                    C@�8��8N�?D             X@)       ,                    :@���Q��?             @*       +                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @.       C                   �T@�ȉo(��??            �V@/       0                    �?Hm_!'1�?#            �H@������������������������       �                     <@1       B                    T@��s����?             5@2       =                    @R���Q�?             4@3       6                   �H@�r����?             .@4       5                    F@�q�q�?             @������������������������       �                      @������������������������       �                     �?7       <                    @I@�8��8��?             (@8       9                   `P@z�G�z�?             @������������������������       �                     @:       ;                   �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @>       ?                    Q@z�G�z�?             @������������������������       �                     @@       A                   @R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     E@E       �                    @K@���b��?v           ��@F       {                    �?8�T����?�            `p@G       Z                   @N@D��T��?\            �`@H       Y                   �I@@4և���?0            �Q@I       J                    @@ףp=
�?$             I@������������������������       �        
             2@K       X                    �J@     ��?             @@L       M                    @F@z�G�z�?             9@������������������������       �                     @N       U                     H@      �?             4@O       T                    @G@      �?              @P       S                    H@r�q��?             @Q       R                    E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @V       W                    E@r�q��?
             (@������������������������       �                      @������������������������       �                     $@������������������������       �                     @������������������������       �                     4@[       \                    @D@X�<ݚ�?,            �O@������������������������       �                     (@]       z                   �Y@��e�B��?%            �I@^       o                   �R@d�
��?!             F@_       n                    �J@�X����?             6@`       e                   �O@���y4F�?             3@a       b                    �G@�q�q�?             @������������������������       �                     �?c       d                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?f       k                    �H@      �?
             0@g       h                   `Q@$�q-�?             *@������������������������       �                     &@i       j                    R@      �?              @������������������������       �                     �?������������������������       �                     �?l       m                   �Q@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @p       w                    @J@���!pc�?             6@q       v                     G@@�0�!��?             1@r       u                   �X@      �?             @s       t                   �T@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     &@x       y                   �S@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @|       �                    @&^�)b�?U             `@}       �                   @K@@�r-��?O            �]@~       �                    �?     ��?
             0@       �                     G@      �?             @������������������������       �                      @�       �                    A@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �E@�q�q�?             (@������������������������       �                     �?�       �                    �J@���!pc�?             &@�       �                    �I@z�G�z�?             $@�       �                   �I@���Q��?             @�       �                   �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �G@l��\��?E            �Y@�       �                    �?�h����?+             L@�       �                   �S@Pa�	�?            �@@�       �                    �E@�����H�?             "@������������������������       �                     @�       �                    R@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     8@������������������������       �                     7@�       �                    V@�㙢�c�?             G@�       �                    �? �q�q�?             8@������������������������       �        	             *@�       �                   �Q@�C��2(�?             &@������������������������       �                      @�       �                     J@�q�q�?             @�       �                   �S@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    @H@�X����?             6@�       �                   `X@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?	             0@�       �                    Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �X@�n_Y�K�?             *@�       �                    �I@z�G�z�?             $@�       �                   `W@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                     H@�eP*L��?             &@�       �                    �C@؇���X�?             @������������������������       �                     @�       �                    W@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       
                   �?�s�n_�?�            �s@�                          `R@��y�S��?w             h@�       �                   �I@dlck+��?t            `g@�       �                     P@,Z0R�?I             ]@�       �                    �N@�ܸb���?;             W@�       �                    @M@D��*�4�?+            @Q@�       �                    �L@�ݜ�?            �C@�       �                   @B@�>����?             ;@�       �                   �?@�<ݚ�?             "@�       �                    8@      �?              @�       �                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �        
             2@�       �                    =@      �?	             (@�       �                    .@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @�       �                    A@�����H�?             "@������������������������       �                     @�       �                   @E@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     >@�       �                    �O@�㙢�c�?             7@�       �                    @O@�S����?             3@�       �                    '@z�G�z�?             @������������������������       �                      @�       �                    >@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    E@؇���X�?             ,@������������������������       �                     (@������������������������       �                      @�       �                    ;@      �?             @������������������������       �                      @�       �                   �A@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@�                          `P@$]��<C�?+            �Q@�       �                   �K@��a�n`�?$             O@�       �                   �J@��
ц��?             *@�       �                     L@�q�q�?             "@������������������������       �                     @�       �                    @O@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �M@      �?             @������������������������       �                     �?������������������������       �                     @�                           P@ZՏ�m|�?            �H@�       �                   �U@��E�B��?            �G@�       �                    @L@������?            �D@�       �                    O@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �M@@-�_ .�?            �B@�       �                    R@�r����?             .@�       �                    @M@�C��2(�?             &@������������������������       �                     "@�       �                   �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �      �?             @������������������������       �                     6@�                         �W@�q�q�?             @�                         �V@�q�q�?             @�                            N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     "@      	                    S@      �?             @                         B@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                         �?j���� �?N            �]@                        �I@����e��?            �@@                         ?@r�q��?             (@������������������������       �                     @                        �D@����X�?             @������������������������       �      �?             @������������������������       �                     @                        �P@؇���X�?             5@������������������������       �                     @                        `R@z�G�z�?             .@                         �L@      �?             @������������������������       �                      @������������������������       �                      @                         �L@�C��2(�?             &@������������������������       �                     @                         @M@r�q��?             @������������������������       �                     �?������������������������       �                     @      :                   @N@��.���?9            �U@      9                   @8�A�0��?             F@      6                   �M@��
ц��?            �C@       +                   �L@4���C�?            �@@!      *                  �T@      �?             2@"      )                  @P@      �?	             (@#      $                   J@և���X�?             @������������������������       �                     @%      (                  @M@      �?             @&      '                   �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @,      1                  @R@�q�q�?             .@-      .                   @M@�<ݚ�?             "@������������������������       �                     @/      0                   I@�q�q�?             @������������������������       �                      @������������������������       �                     @2      3                  `U@      �?             @������������������������       �                     �?4      5                  �W@���Q��?             @������������������������       �      �?             @������������������������       �                     �?7      8                  �P@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @;      @                   �N@0,Tg��?             E@<      ?                   @�8��8��?             (@=      >                   L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @A      N                  @N@�q�q�?             >@B      M                   @���y4F�?             3@C      J                    R@������?             1@D      I                   �P@؇���X�?
             ,@E      F                  �9@      �?              @������������������������       �                     �?G      H                    P@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @K      L                  �?@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @O      T                    P@�eP*L��?	             &@P      Q                  �T@����X�?             @������������������������       �                     @R      S                   �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @U      X                   @      �?             @V      W                   S@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?q�tq�bh�h"h#K �q�h%�q�Rq�(KMYKK�q�hV�B�        t@     �y@     @[@     �I@      4@      F@      0@      F@      (@      &@      (@      "@      @      @      @              �?      @              @      �?      @      �?       @               @       @       @              �?       @      �?      @              @      �?      @                      �?               @      @     �@@      @       @       @       @              @       @      @      �?      @      �?                      @      �?              �?              �?      9@              *@      �?      (@              @      �?      @      �?                      @      @             @V@      @       @      @       @      �?       @                      �?               @     �U@      @     �F@      @      <@              1@      @      1@      @      *@       @       @      �?       @                      �?      &@      �?      @      �?      @              �?      �?              �?      �?              @              @      �?      @              �?      �?              �?      �?                      �?      E@             �j@     �v@     @a@      _@     �@@      Y@      @     @P@      @     �F@              2@      @      ;@      @      4@              @      @      .@      @      @      �?      @      �?      �?              �?      �?                      @       @               @      $@       @                      $@              @              4@      <@     �A@              (@      <@      7@      5@      7@      .@      @      .@      @      �?       @              �?      �?      �?      �?                      �?      ,@       @      (@      �?      &@              �?      �?              �?      �?               @      �?      �?      �?      �?                      @      @      0@      @      ,@      @      @      @      �?              �?      @                       @              &@      @       @               @      @              @             @Z@      8@      Y@      2@      @      "@      @      �?       @              �?      �?              �?      �?              @       @      �?              @       @       @       @       @      @       @      �?              �?       @                       @              @      �?             @W@      "@     �K@      �?      @@      �?       @      �?      @               @      �?       @                      �?      8@              7@              C@       @      7@      �?      *@              $@      �?       @               @      �?      �?      �?              �?      �?              �?              .@      @      @      �?              �?      @              $@      @       @      �?       @                      �?       @      @       @       @      @       @               @      @              @                      @      @      @      �?      @              @      �?      @              @      �?              @             �R@     �m@      :@     �d@      7@     �d@      "@     �Z@      "@     �T@      @      P@      @      A@       @      9@       @      @      �?      @      �?       @               @      �?                      @      �?                      2@      @      "@       @      �?      �?              �?      �?      �?       @              @      �?      @      �?       @               @              >@      @      3@      @      0@      �?      @               @      �?       @      �?                       @       @      (@              (@       @              �?      @               @      �?      �?      �?                      �?              8@      ,@     �L@      ,@      H@      @      @      @      @              @      @       @      @                       @      @      �?              �?      @               @     �D@      @     �D@      @     �B@       @       @               @       @               @     �A@       @      *@      �?      $@              "@      �?      �?      �?                      �?      �?      @              6@       @      @       @      �?      �?      �?      �?                      �?      �?                      @       @                      "@      @      @      @      �?              �?      @                       @     �H@     �Q@      4@      *@       @      $@              @       @      @       @       @              @      2@      @      @              (@      @       @       @               @       @              $@      �?      @              @      �?              �?      @              =@     �L@      2@      :@      2@      5@      ,@      3@      "@      "@      @      "@      @      @              @      @      �?      �?      �?              �?      �?               @                      @      @              @      $@       @      @              @       @      @       @                      @      @      @      �?               @      @       @       @              �?      @       @      @                       @              @      &@      ?@      �?      &@      �?      @              @      �?                      @      $@      4@      @      .@      @      *@       @      (@       @      @      �?              �?      @              @      �?                      @       @      �?              �?       @                       @      @      @      @       @      @              �?       @      �?                       @      �?      @      �?       @               @      �?                      �?q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       r   tr  bK�r  Rr  }r  (hKhjM�hkh"h#K �r  h%�r  Rr  (KM��r  hr�BU         �                    �?4�5����?�           ��@       3                    �?����&�?           Py@                            K@f���M�?*             O@                            E@�G��l��?             5@������������������������       �                     @                          �M@ҳ�wY;�?             1@                          �<@      �?             $@������������������������       �                      @	       
                     G@      �?              @������������������������       �                     �?                          �A@����X�?             @������������������������       �                     @                          @F@      �?             @                           �H@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     �?                           �I@؇���X�?             @                           @H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @       2                    �P@���� �?            �D@       #                   �S@�θ�?            �C@       "                   �N@      �?             8@       !                   @L@�θ�?             *@                          @F@�C��2(�?             &@������������������������       �                     @                            N@r�q��?             @������������������������       �                     @                           �G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@$       1                   �V@���Q��?
             .@%       0                    �O@�eP*L��?             &@&       /                    V@X�<ݚ�?             "@'       (                    @M@����X�?             @������������������������       �                     �?)       .                    U@r�q��?             @*       +                   `T@�q�q�?             @������������������������       �                     �?,       -                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @4       o                    �I@��qqI��?�            pu@5       :                    @C@y�w[��?C            @[@6       7                    @B@@4և���?
             ,@������������������������       �                     @8       9                    �B@؇���X�?             @������������������������       �                     �?������������������������       �                     @;       ^                    �G@��̅��?9            �W@<       O                   @P@F�����?"            �L@=       @                    �D@l��
I��?             ;@>       ?                   @I@�q�q�?             @������������������������       �                      @������������������������       �                     �?A       F                   �G@      �?             8@B       C                   @E@���Q��?             $@������������������������       �                      @D       E                    @F@      �?              @������������������������       �                     @������������������������       �                     @G       L                    @G@؇���X�?	             ,@H       I                    J@�8��8��?             (@������������������������       �                     @J       K                    @F@z�G�z�?             @������������������������       �                     �?������������������������       �                     @M       N                   @I@      �?              @������������������������       �                     �?������������������������       �                     �?P       U                   �Q@���Q��?             >@Q       R                     E@      �?             (@������������������������       �                     @S       T                    @F@և���X�?             @������������������������       �                     @������������������������       �                     @V       W                    �D@      �?             2@������������������������       �                     @X       Y                    �E@�	j*D�?	             *@������������������������       �                     @Z       [                    @F@�q�q�?             @������������������������       �                     @\       ]                   `R@�q�q�?             @������������������������       �                     �?������������������������       �                      @_       b                    @H@�d�����?             C@`       a                   �X@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @c       d                   �K@`�Q��?             9@������������������������       �                     &@e       f                    P@և���X�?	             ,@������������������������       �                     @g       l                    @I@�q�q�?             "@h       i                   `P@���Q��?             @������������������������       �                      @j       k                   �Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?m       n                   @Z@      �?             @������������������������       �                     @������������������������       �                     �?p       �                    R@��O
�?�            @m@q       t                    @(�Y7B��?�            `i@r       s                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @u       �                   �I@      �?�             i@v       �                   @F@���	���?Z             a@w       �                    �R@t����?F            �Z@x       �                   �E@ȵHPS!�?D             Z@y       z                    +@ i���t�?@            �X@������������������������       �        
             .@{       �                    .@�gc� �?6            �T@|       }                    �N@      �?             @������������������������       �                     �?~                           @O@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @C@$��$�L�?3            �S@�       �                    @M@<���D�?+            �P@�       �                    @L@��G���?            �B@�       �                    @J@      �?             8@������������������������       �                     @�       �                   �A@R���Q�?             4@������������������������       �                     ,@�       �                   �B@      �?             @�       �                   @B@���Q��?             @�       �                    @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    �L@�	j*D�?	             *@�       �                    8@      �?             @�       �                   �3@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �@@؇���X�?             @������������������������       �                      @�       �                   @B@z�G�z�?             @������������������������       �      �?             @������������������������       �                     �?�       �                   @@@XB���?             =@�       �                   �>@      �?
             0@������������������������       �                     $@�       �                    �O@r�q��?             @������������������������       �                     @�       �                     P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             *@������������������������       �                     *@�       �                    @M@�q�q�?             @������������������������       �                     @������������������������       ��q�q�?             @�       �                    B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ?@�       �                   @K@��s����?+            �O@�       �                   �J@���Q��?             $@�       �                    @L@�q�q�?             @������������������������       �                     @�       �                   @J@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �O@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �P@f1r��g�?#            �J@�       �                     P@��s����?             E@�       �                    @L@�ݜ�?            �C@�       �                    @K@      �?
             (@�       �                   @N@�����H�?             "@�       �                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    O@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @M@�>����?             ;@������������������������       �                     "@�       �                   �N@�����H�?             2@�       �                    �N@���Q��?             @�       �                    �M@�q�q�?             @������������������������       �                     �?�       �                   �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     @������������������������       �                     &@�       �                   `R@�4�����?             ?@�       �                    �L@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �Y@������?             ;@�       �                   �R@�θ�?             :@������������������������       �                     @�       �                    �M@�z�G��?             4@�       �                    U@�eP*L��?             &@�       �                   @T@      �?              @�       �                    �J@      �?             @������������������������       �                      @�       �                    �K@      �?             @������������������������       �                      @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     �?�       �       
             �?������?�            �t@�       �                     R@�FVQ&�?=            �X@�       �                    �G@h�a��?;            @X@������������������������       �                     B@�       �                    �H@85�}C�?&            �N@�       �                   @U@����X�?             @�       �                   �Q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    C@�X�<ݺ?"             K@�       �                   �7@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                    �H@�       �                    `R@      �?              @������������������������       �                     �?������������������������       �                     �?�                          �J@ڷv���?�            �l@�                          @K@      �?(             L@�       �                    A@�����?             3@������������������������       �                     @�       �                    �?և���X�?             ,@������������������������       �                     @�       �                    �G@�q�q�?             "@������������������������       �                     �?�       �                   @F@      �?              @������������������������       �                     @�                          �I@�q�q�?             @������������������������       �                      @������������������������       �                     �?                         @���@��?            �B@                        �E@r֛w���?             ?@                         �Q@j���� �?             1@                         �L@����X�?             ,@������������������������       �                     �?                          N@�θ�?             *@                         �?���Q��?             @	      
                   ?@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @                         @M@      �?              @������������������������       �                     �?������������������������       �                     �?                         �?      �?              @������������������������       �                      @                         @O@r�q��?             @                         $@�q�q�?             @������������������������       �                     �?                         �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @                        �G@@4և���?             ,@                         @N@      �?              @                        �F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @!      d                   �K@����S��?v            �e@"      3                   �F@     �?V             `@#      0                   @pH����?+            �P@$      '                  �P@     p�?(             P@%      &                  @P@���!pc�?             &@������������������������       �                      @������������������������       �                     @(      /                  �U@�&=�w��?!            �J@)      *                  �T@�C��2(�?             6@������������������������       �        	             0@+      .                   @C@�q�q�?             @,      -                   @@@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     ?@1      2                   �C@�q�q�?             @������������������������       �                      @������������������������       �                     �?4      M                   �I@�̚��?+            �N@5      :                  �S@�f7�z�?             =@6      9                   @r�q��?             @7      8                  �Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @;      H                   �H@8����?             7@<      G                   @������?             1@=      @                  �W@     ��?
             0@>      ?                   W@���Q��?             @������������������������       �                     @������������������������       �                      @A      B                   @H@�C��2(�?             &@������������������������       �                     @C      D                   �?      �?             @������������������������       �                     �?E      F                  �X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?I      L                   @I@      �?             @J      K                   �?���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     �?N      c                   @     ��?             @@O      T                   �J@V�a�� �?             =@P      Q                   �?$�q-�?
             *@������������������������       �                     @R      S                  @Y@؇���X�?             @������������������������       �                     @������������������������       �                     �?U      \                   �?     ��?             0@V      Y                   @K@�q�q�?             "@W      X                   W@���Q��?             @������������������������       �                     @������������������������       �                      @Z      [                   R@      �?             @������������������������       �                     �?������������������������       �                     @]      b                  @S@����X�?             @^      _                  @M@�q�q�?             @������������������������       �                     �?`      a                   @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @e      n                   �?\X��t�?              G@f      g                   �L@�θ�?             *@������������������������       �                     @h      i                  @L@�q�q�?             "@������������������������       �                     �?j      m                   @M@      �?              @k      l                  @T@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @o      p                  �L@:ɨ��?            �@@������������������������       �                     @q      �                   @V�a�� �?             =@r      w                   S@��s����?             5@s      v                   P@�C��2(�?             &@t      u                  �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@x      y                   �L@�z�G��?             $@������������������������       �                     �?z                         �P@�<ݚ�?             "@{      |                   �N@      �?              @������������������������       �                     @}      ~                   �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                   �O@      �?              @������������������������       �                     @�      �                  �V@�q�q�?             @������������������������       �                      @������������������������       �                     �?r	  tr
  bh�h"h#K �r  h%�r  Rr  (KM�KK�r  hV�BP       �t@     y@      X@     Ps@      6@      D@      &@      $@              @      &@      @      @      @       @              @      @      �?               @      @              @       @       @       @      �?      �?              �?      �?              �?      @      �?       @      �?       @                      �?      @              &@      >@      "@      >@      @      5@      @      $@      �?      $@              @      �?      @              @      �?      �?      �?                      �?       @                      &@      @      "@      @      @      @      @       @      @      �?              �?      @      �?       @              �?      �?      �?              �?      �?                      @       @               @                      @       @             �R@     �p@     �B@      R@      �?      *@              @      �?      @      �?                      @      B@     �M@      :@      ?@       @      3@       @      �?       @                      �?      @      2@      @      @               @      @      @              @      @               @      (@      �?      &@              @      �?      @      �?                      @      �?      �?              �?      �?              2@      (@      "@      @      @              @      @              @      @              "@      "@              @      "@      @      @               @      @              @       @      �?              �?       @              $@      <@       @      &@              &@       @               @      1@              &@       @      @      @              @      @       @      @               @       @      �?       @                      �?      �?      @              @      �?             �B@     �h@      ;@      f@       @      �?              �?       @              9@     �e@      *@      _@      *@     @W@      (@      W@      $@      V@              .@      $@     @R@       @       @              �?       @      �?       @                      �?       @     �Q@       @      M@      @      >@      @      5@              @      @      1@              ,@      @      @       @      @       @      �?              �?       @                       @      �?              @      "@      @      @      @      �?              �?      @                       @      �?      @               @      �?      @      �?      @              �?      �?      <@      �?      .@              $@      �?      @              @      �?       @      �?                       @              *@              *@       @      @              @       @      �?      �?      �?              �?      �?                      ?@      (@     �I@      @      @       @      @              @       @      �?       @                      �?       @       @               @       @               @     �F@       @      A@      @      A@      @      "@      �?       @      �?       @               @      �?                      @       @      �?              �?       @               @      9@              "@       @      0@       @      @       @      �?      �?              �?      �?              �?      �?                       @              *@      @                      &@      $@      5@      @      �?      @                      �?      @      4@      @      4@              @      @      ,@      @      @      @      @      @      @               @      @      �?       @              �?      �?              �?      �?                       @      @                      "@      �?             �m@      W@     @W@      @      W@      @      B@              L@      @      @       @       @       @       @                       @      @             �I@      @       @      @       @                      @     �H@              �?      �?              �?      �?              b@     �U@      5@     �A@      *@      @      @               @      @      @              @      @      �?               @      @              @       @      �?       @                      �?       @      =@       @      7@      @      $@      @      $@      �?              @      $@       @      @      �?       @              �?      �?      �?      �?      �?              �?      �?              �?      @               @      �?      @      �?       @              �?      �?      �?              �?      �?                      @      @              �?      *@      �?      @      �?      �?              �?      �?                      @              @              @     �^@     �I@     �Y@      9@      N@      @     �M@      @       @      @       @                      @     �I@       @      4@       @      0@              @       @      �?       @      �?                       @      @              ?@              �?       @               @      �?             �E@      2@      1@      (@      �?      @      �?       @      �?                       @              @      0@      @      *@      @      *@      @      @       @      @                       @      $@      �?      @              @      �?      �?               @      �?       @                      �?              �?      @      @       @      @      �?              �?      @      �?              :@      @      7@      @      (@      �?      @              @      �?      @                      �?      &@      @      @      @      @       @      @                       @      @      �?              �?      @              @       @      �?       @              �?      �?      �?              �?      �?              @              @              4@      :@      $@      @      @              @      @              �?      @       @      �?       @      �?                       @      @              $@      7@      @              @      7@      @      1@      �?      $@      �?      �?              �?      �?                      "@      @      @      �?               @      @      �?      @              @      �?       @      �?                       @      �?               @      @              @       @      �?       @                      �?r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h<Kh=Kh>h"h#K �r  h%�r  Rr  (KK�r  hV�C              �?r  tr  bhJhZhEC       r  �r  Rr  h^Kh_h`Kh"h#K �r  h%�r  Rr  (KK�r  hE�C       r   tr!  bK�r"  Rr#  }r$  (hKhjMUhkh"h#K �r%  h%�r&  Rr'  (KMU�r(  hr�B�J         �                   @L@6������?�           ��@                           �?ƆQ����?�            s@                           C@H�z�G�?             D@       	                    �?�q�q�?             (@                           5@�q�q�?             "@������������������������       �                      @                          �A@؇���X�?             @������������������������       �                     @������������������������       ��q�q�?             @
                          �7@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?��X��?             <@                           J@�eP*L��?             &@                           E@z�G�z�?             @������������������������       �                      @                            M@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �H@r�q��?             @                            F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?@�0�!��?             1@������������������������       �                     @                          @G@�z�G��?             $@������������������������       �                     @                           �O@      �?             @������������������������       �                     �?������������������������       �                     @        g                    �?�	M���?�            �p@!       V                   �I@°	~��?{             h@"       %                     E@�}#���?j            �d@#       $                   �D@      �?              @������������������������       �                     �?������������������������       �                     �?&       )                    @���C"��?h            �d@'       (                    @���Q��?             @������������������������       �                     @������������������������       �                      @*       +                    @J@D���D|�?e            �c@������������������������       �                     =@,       /                    �J@��a�!��?R            @`@-       .                    E@���Q��?             @������������������������       �                     @������������������������       �                      @0       1                    *@H�̱���?O            @_@������������������������       �                     0@2       3                    @L@p���h�?I            @[@������������������������       �                     ?@4       U                     P@��-�=��?7            �S@5       F                    �N@(2��R�?*            �M@6       A                    @M@ףp=
�?             >@7       <                    �L@      �?             0@8       ;                   @@@ףp=
�?             $@9       :                    :@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @=       >                   �@@r�q��?             @������������������������       �                     @?       @                   @B@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?B       C                   �E@@4և���?             ,@������������������������       �                     "@D       E                   �F@z�G�z�?             @������������������������       �      �?              @������������������������       �                     @G       P                    �O@д>��C�?             =@H       I                    .@z�G�z�?             4@������������������������       �                      @J       K                   �E@�����H�?             2@������������������������       �                     *@L       M                    @O@���Q��?             @������������������������       �                      @N       O                   @G@�q�q�?             @������������������������       �                      @������������������������       �                     �?Q       R                   �=@�����H�?             "@������������������������       �                     @S       T                   �?@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@W       b                   �K@�5��?             ;@X       [                   @J@���Q��?             .@Y       Z                    �J@      �?             @������������������������       �                      @������������������������       �                      @\       a                    �M@���|���?             &@]       `                   �J@և���X�?             @^       _                    �H@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @c       d                    �G@r�q��?	             (@������������������������       �                     @e       f                    @K@����X�?             @������������������������       �                      @������������������������       �                     @h       q                    �?<ݚ)�?&             R@i       j                   �8@և���X�?             5@������������������������       �                     @k       p                     P@      �?
             0@l       o                   @@@$�q-�?             *@m       n                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     @r       �                    @��x_F-�?            �I@s       ~                   �E@z�G�z�?            �F@t       }                   �D@�LQ�1	�?             7@u       v                    �N@      �?
             4@������������������������       �                     @w       |                   �C@X�Cc�?             ,@x       {                   �1@      �?             (@y       z                    $@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @       �                   �G@���7�?             6@�       �                     P@ףp=
�?             $@������������������������       �                     @�       �                   �F@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@�       �                    �K@r�q��?             @������������������������       �                     �?������������������������       �                     @�                           @L@��V�9�?           �z@�       �                    �?0e­���?�            pr@�       �                    @C@���H��?5             U@�       �                    �?���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                    T@�L���?.            �R@�       �                   �S@6YE�t�?            �@@�       �                   �P@      �?             @@������������������������       �                     "@�       �                    �?�㙢�c�?             7@�       �                   @Q@z�G�z�?             @������������������������       �                      @�       �                   @R@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             2@������������������������       �                     �?�       �                    �?��Y��]�?            �D@������������������������       �                     9@�       �                   �W@      �?
             0@������������������������       �                     $@�       �                   @X@r�q��?             @�       �                    @I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�V�K���?�            `j@�       �                   �R@�G�z�?0             T@�       �                    @F@�G�z��?             D@�       �                    �C@�C��2(�?             &@�       �                   �O@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                      @�       �                   `P@�f7�z�?             =@�       �                    �H@���!pc�?             &@������������������������       �                     �?�       �                   �O@z�G�z�?             $@�       �                   �M@      �?              @������������������������       �                     �?�       �                   @N@����X�?             @�       �                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �I@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �J@�<ݚ�?             2@�       �                    @H@@4և���?             ,@������������������������       �                     @�       �                    �I@      �?              @������������������������       �z�G�z�?             @������������������������       �                     @�       �                   �P@      �?             @�       �                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                     E@z�G�z�?             D@�       �                   @W@P���Q�?             4@������������������������       �        	             1@�       �                    @C@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �E@��Q��?             4@������������������������       �                     @�       �                    Z@������?
             1@�       �                    T@�r����?             .@������������������������       �                     "@�       �                   `T@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    @F@�������?U            ``@�       �                    �? 7���B�?$             K@�       �                    �B@�FVQ&�?            �@@�       �                   �V@8�Z$���?             *@�       �                   �T@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     4@������������������������       �                     5@�       �                    �H@��مD�?1            @S@�       �                    @      �?             8@�       �                   �X@���Q��?             4@�       �                    @G@����X�?
             ,@�       �                   �R@      �?              @�       �                    Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �W@      �?             @�       �                    �?      �?             @������������������������       �                      @�       �                   �Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @H@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?0��_��?!            �J@������������������������       �                     =@�       �                    @�q�q�?             8@�       �                    @K@z�G�z�?             4@�       �                   �X@��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?�       �                   @P@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �K@      �?             @�       �                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                        �L@|��Q��?V            �`@������������������������       �                     @                         �?�lg����?S             `@                         �?      �?             @@                        �V@���|���?             6@                         `P@D�n�3�?             3@                         V@ҳ�wY;�?             1@      	                   �O@8�Z$���?	             *@������������������������       �                      @
                        �R@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @                        @R@z�G�z�?             $@                         �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @      0                   �?�Y �K�??            @X@                        @P@r�q��?             H@                        @M@�q�q�?             "@������������������������       �                     @                        �N@      �?             @������������������������       �                     �?                          P@���Q��?             @������������������������       �                     @������������������������       �                      @      /                  �W@�ݜ�?            �C@      (                   �M@     ��?             @@       #                    M@���|���?             &@!      "                   U@z�G�z�?             @������������������������       �                     @������������������������       �                     �?$      '                   U@      �?             @%      &                  @R@���Q��?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     �?)      *                    P@���N8�?             5@������������������������       �        
             ,@+      .                   `P@؇���X�?             @,      -                  �R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @1      8                   �?�`���?             �H@2      7                   @M@����X�?	             ,@3      6                   �L@z�G�z�?             @4      5                  �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@9      J                   @N@���Q��?            �A@:      =                  �P@�X����?             6@;      <                   �M@�q�q�?             @������������������������       �                     �?������������������������       �                      @>      I                   �M@�d�����?             3@?      B                   U@     ��?	             0@@      A                    M@�q�q�?             @������������������������       �                     �?������������������������       �                      @C      H                   @M@�θ�?             *@D      E                   V@      �?              @������������������������       �                     �?F      G                  �W@����X�?             @������������������������       ����Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @K      T                    Q@��
ц��?
             *@L      M                  @N@�q�q�?	             (@������������������������       �                     @N      Q                   @�<ݚ�?             "@O      P                   T@r�q��?             @������������������������       �                     @������������������������       �                     �?R      S                  �Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?r)  tr*  bh�h"h#K �r+  h%�r,  Rr-  (KMUKK�r.  hV�BP       �t@     �x@     �Q@     `m@      7@      1@      @       @      @      @       @              �?      @              @      �?       @      �?       @      �?                       @      3@      "@      @      @      @      �?       @               @      �?              �?       @              �?      @      �?      �?              �?      �?                      @      ,@      @      @              @      @      @              �?      @      �?                      @     �G@     @k@      9@      e@      ,@      c@      �?      �?      �?                      �?      *@     �b@       @      @              @       @              &@     �b@              =@      &@     �]@      @       @      @                       @       @     @]@              0@       @     @Y@              ?@       @     �Q@       @     �I@      @      ;@       @      ,@      �?      "@      �?      @              @      �?                      @      �?      @              @      �?       @      �?      �?              �?      �?      *@              "@      �?      @      �?      �?              @      @      8@      @      0@       @               @      0@              *@       @      @               @       @      �?       @                      �?      �?       @              @      �?      @      �?                      @              3@      &@      0@      "@      @       @       @               @       @              @      @      @      @      @      �?      @                      �?              @      @               @      $@              @       @      @       @                      @      6@      I@      (@      "@              @      (@      @      (@      �?       @      �?       @                      �?      $@                      @      $@     �D@      "@      B@       @      .@      @      .@              @      @      "@      @      "@      @      �?              �?      @                       @       @              @              �?      5@      �?      "@              @      �?      @              @      �?                      (@      �?      @      �?                      @     �p@     �d@     �j@     �T@     �R@      $@      @      @              @      @              Q@      @      <@      @      <@      @      "@              3@      @      �?      @               @      �?       @      �?                       @      2@                      �?      D@      �?      9@              .@      �?      $@              @      �?       @      �?              �?       @              @             @a@     @R@      :@      K@      2@      6@      �?      $@      �?       @              �?      �?      �?               @      1@      (@      @       @      �?               @       @       @      @              �?       @      @      �?       @               @      �?              �?      @      �?                      @               @      ,@      @      *@      �?      @              @      �?      @      �?      @              �?      @      �?       @               @      �?                      �?       @      @@      �?      3@              1@      �?       @      �?                       @      @      *@      @              @      *@       @      *@              "@       @      @       @                      @       @              \@      3@      J@       @      ?@       @      &@       @      �?       @      �?                       @      $@              4@              5@              N@      1@      (@      (@      (@       @      $@      @      @      �?       @      �?       @                      �?      @              @      @      �?      @               @      �?      �?      �?                      �?       @               @      @       @                      @              @      H@      @      =@              3@      @      0@      @      ,@      �?      ,@                      �?       @      @       @                      @      @      �?      �?      �?      �?                      �?       @             �J@     @T@      @              H@     @T@      0@      0@       @      ,@       @      &@      @      &@       @      &@               @       @      @              @       @              @               @                      @       @       @      �?       @               @      �?              @              @@     @P@       @      D@      @      @              @      @      @      �?               @      @              @       @              @      A@      @      ;@      @      @      �?      @              @      �?              @      @      @       @      �?       @       @                      �?      �?      4@              ,@      �?      @      �?      �?      �?                      �?              @              @      8@      9@      $@      @      �?      @      �?      �?      �?                      �?              @      "@              ,@      5@      @      .@       @      �?              �?       @              @      ,@      @      &@       @      �?              �?       @              @      $@      @      @      �?               @      @       @      @               @              @              @      @      @      @      @              @      @       @      @      �?      @                      �?       @      �?       @                      �?              �?r/  tr0  bubhhubh)�r1  }r2  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h<Kh=Kh>h"h#K �r3  h%�r4  Rr5  (KK�r6  hV�C              �?r7  tr8  bhJhZhEC       r9  �r:  Rr;  h^Kh_h`Kh"h#K �r<  h%�r=  Rr>  (KK�r?  hE�C       r@  trA  bK�rB  RrC  }rD  (hKhjM?hkh"h#K �rE  h%�rF  RrG  (KM?�rH  hr�B�E         �                    �?U�ք�?�           ��@                           �?r=ά�{�?�            Px@                          @L@�q�q�?&             N@                           ;@r�q��?             8@������������������������       �                      @                           @I@�C��2(�?             6@                          �A@�<ݚ�?             "@������������������������       �                      @	                          @H@����X�?             @
                          @C@���Q��?             @������������������������       �      �?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@                           @M@�q�q�?             B@                          �T@      �?             8@                          �Q@և���X�?
             ,@������������������������       �                     @                           @H@؇���X�?             @                            E@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@                           S@      �?             (@������������������������       �                     @                           �N@�q�q�?             "@������������������������       �                     @                           @P@      �?             @������������������������       �                     @������������������������       �                     @        M                   @J@��^�V��?�            �t@!       "                   �:@�f"Nf�?l             f@������������������������       �                    �D@#       L                    �R@�IєX�?T             a@$       3                    �G@X�Հ�+�?S            �`@%       &                    @D@�����H�?             ;@������������������������       �                     "@'       (                    �D@r�q��?             2@������������������������       �                     �?)       0                    @G@�t����?
             1@*       /                    H@@4և���?             ,@+       ,                    E@      �?              @������������������������       �                     @-       .                    @F@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @1       2                   @I@�q�q�?             @������������������������       �                      @������������������������       �                     �?4       5                    @L@ 7���B�?D             [@������������������������       �                     D@6       ;                    �L@�IєX�?-             Q@7       8                    A@�q�q�?             @������������������������       �                     �?9       :                    H@z�G�z�?             @������������������������       �                     @������������������������       �                     �?<       =                    @O@�g�y��?)             O@������������������������       �                     <@>       G                    F@�IєX�?             A@?       F                   @@@(;L]n�?             >@@       A                   �>@�����H�?             "@������������������������       �                     @B       E                     P@      �?             @C       D                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     5@H       K                   @G@      �?             @I       J                     P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?N       Y                    �D@���=A�?a             c@O       P                     B@$�q-�?             :@������������������������       �                     "@Q       R                    �B@�t����?             1@������������������������       �                     �?S       X                    Q@      �?             0@T       U                    @C@z�G�z�?             @������������������������       �                      @V       W                   @P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             &@Z       �                   �Y@�ՙ/�?N            �_@[       �                    `P@P&��?H            �]@\       �                   �R@r���@�?A            �Z@]       ^                   �J@^|�_��?,            �Q@������������������������       �                      @_       �                    R@������?+            @Q@`       �                   �P@*;L]n�?&             N@a       b                    �F@Np�����?            �I@������������������������       �                     @c       d                    �G@�q���?             H@������������������������       �                     @e       �                   �P@�ݏ^���?            �F@f                          `P@��6���?             E@g       z                   @O@���>4��?             <@h       s                    �M@�G��l��?             5@i       j                   �K@      �?             (@������������������������       �                     @k       n                   @M@�q�q�?             "@l       m                     M@      �?              @������������������������       �                     �?������������������������       �                     �?o       p                   @N@����X�?             @������������������������       �                      @q       r                    �I@���Q��?             @������������������������       �                      @������������������������       �                     @t       u                    �N@�<ݚ�?             "@������������������������       �                     @v       y                   �K@���Q��?             @w       x                    �O@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?{       ~                    P@����X�?             @|       }                     L@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                    @K@����X�?             ,@������������������������       �                     @�       �                    �M@      �?              @������������������������       �                     @�       �                     P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @I@�����H�?             "@�       �                    �F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   `R@�q�q�?             "@�       �                    @H@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �L@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �W@tk~X��?             B@�       �                    @J@��a�n`�?             ?@�       �                   �U@�IєX�?             1@������������������������       �                     *@�       �                    V@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �K@և���X�?
             ,@������������������������       �                     @�       �                   �V@z�G�z�?             $@�       �                    �M@�����H�?             "@�       �                    �L@      �?             @������������������������       �                     �?�       �                   �U@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                     K@      �?              @������������������������       �                     @������������������������       �                     �?�       �                   �J@ �>�?�            �u@�       �                    �?�D����?5             U@�       �                    @�θ�?             :@�       �                   @C@���!pc�?             6@�       �                    �M@؇���X�?             @������������������������       �                     @�       �                   �7@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@������������������������       �                     @�       �                     K@>���Rp�?&             M@�       �                   @I@     ��?             0@�       �                    A@������?             .@������������������������       �                     @�       �                   �D@�q�q�?	             (@������������������������       �                      @�       �                   �E@z�G�z�?             $@������������������������       �                      @�       �                    �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                    �?@4և���?             E@������������������������       �                     "@�       �                   �G@�C��2(�?            �@@�       �                   �F@      �?             8@�       �                    @�C��2(�?             6@�       �                     N@ףp=
�?             4@������������������������       �                     �?�       �                    D@�}�+r��?
             3@������������������������       �                     (@�       �                   �E@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �       	             �?D�~�.��?�            Pp@�       �                   @X@������?2            �T@�       �                   �W@`Jj��?'             O@�       �                     N@XB���?$             M@�       �                    �?p���?             I@������������������������       �                     @@�       �                    �H@�X�<ݺ?             2@������������������������       �                     "@�       �                    @I@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                    @      �?              @������������������������       �                     @������������������������       �                     �?�       �                     G@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     4@�       ,                  �X@؀2��a�?s            `f@�                          �?�ګH9�?]            �a@�       �                   �K@\#r��?)            �N@������������������������       �                     �?�                         �W@�8��8��?(             N@�       �                    W@ i���t�?             �H@�       �                   �U@dP-���?            �G@�       �                   �T@��-�=��?            �C@�       �                   �P@`Jj��?             ?@�       �                     C@�����H�?             2@������������������������       �                     �?�       �                    @L@�IєX�?
             1@������������������������       �                     $@�       �                    �M@؇���X�?             @�       �                   �P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �        	             *@�       �                     K@      �?              @�       �                    �B@؇���X�?             @�       �                    @@@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @                          �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@      !                   @��}*_��?4            @T@      
                   P@L
�q��?'            �M@                         �L@@4և���?             ,@������������������������       �                     $@      	                  @N@      �?             @������������������������       �                     �?������������������������       �                     @                         S@k��9�?            �F@                         �E@�d�����?             3@������������������������       �                     �?                         �M@�<ݚ�?
             2@������������������������       �                      @                         @P@���Q��?             $@                         �N@z�G�z�?             @                        �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         �V@���B���?             :@                        �U@�E��ӭ�?             2@                          I@     ��?
             0@                         @F@�q�q�?             "@������������������������       �                     @                         T@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @"      '                  �Q@�eP*L��?             6@#      &                  @O@����X�?             ,@$      %                   �O@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @(      )                   @J@      �?              @������������������������       �                     @*      +                   �L@���Q��?             @������������������������       �                      @������������������������       �                     @-      6                    H@��J�fj�?            �B@.      1                   @A@      �?             4@/      0                  �Z@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @2      5                  �Y@�C��2(�?	             &@3      4                   Y@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @7      :                   �?ҳ�wY;�?             1@8      9                  �[@      �?              @������������������������       �                     @������������������������       �                     @;      >                   Y@�����H�?             "@<      =                   @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @rI  trJ  bh�h"h#K �rK  h%�rL  RrM  (KM?KK�rN  hV�B�        t@     �y@     �T@      s@      9@     �A@      @      4@       @               @      4@       @      @               @       @      @       @      @      �?      @      �?                       @              *@      5@      .@      2@      @       @      @      @              �?      @      �?       @               @      �?                      @      $@              @      "@              @      @      @              @      @      @      @                      @      M@     �p@       @      e@             �D@       @      `@      @      `@      @      8@              "@      @      .@      �?               @      .@      �?      *@      �?      @              @      �?      @              @      �?                      @      �?       @               @      �?              @      Z@              D@      @      P@       @      @      �?              �?      @              @      �?               @      N@              <@       @      @@      �?      =@      �?       @              @      �?      @      �?      �?              �?      �?                       @              5@      �?      @      �?       @      �?                       @              �?      �?              I@     �Y@       @      8@              "@       @      .@      �?              �?      .@      �?      @               @      �?       @               @      �?                      &@      H@     �S@     �D@     @S@     �D@     �P@      A@     �B@       @              @@     �B@      :@      A@      9@      :@              @      9@      7@      @              6@      7@      3@      7@      .@      *@      $@      &@      @      "@              @      @      @      �?      �?              �?      �?               @      @               @       @      @       @                      @      @       @      @              @       @      @      �?              �?      @                      �?      @       @      @       @      @                       @      �?              @      $@              @      @      @      @              �?      @              @      �?              @              �?       @      �?       @               @      �?                      @      @      @      @      �?              �?      @               @       @       @                       @      @      =@      @      8@      �?      0@              *@      �?      @      �?                      @      @       @      @               @       @      �?       @      �?      @              �?      �?       @      �?                       @              @      �?                      @              &@      @      �?      @                      �?     �m@     �Z@      A@      I@      4@      @      0@      @      �?      @              @      �?       @      �?                       @      .@              @              ,@      F@      &@      @      &@      @      @               @      @               @       @       @       @              @       @      @                       @              �?      @     �C@              "@      @      >@      @      5@       @      4@       @      2@      �?              �?      2@              (@      �?      @      �?                      @               @      �?      �?      �?                      �?              "@     �i@      L@     �S@      @      M@      @      L@       @     �H@      �?      @@              1@      �?      "@               @      �?              �?       @              @      �?      @                      �?       @       @       @                       @      4@             �_@      J@     �Z@      B@     �K@      @              �?     �K@      @      F@      @     �E@      @     �A@      @      =@       @      0@       @              �?      0@      �?      $@              @      �?      @      �?      @                      �?       @              *@              @       @      @      �?       @      �?       @                      �?      @                      �?       @              �?      �?      �?                      �?      &@             �I@      >@     �C@      4@      *@      �?      $@              @      �?              �?      @              :@      3@      @      ,@      �?              @      ,@               @      @      @      @      �?      �?      �?      �?                      �?      @                      @      5@      @      *@      @      *@      @      @      @      @              �?      @              @      �?              @                       @       @              (@      $@      $@      @      @      @              @      @              @               @      @              @       @      @       @                      @      5@      0@      .@      @      @      @              @      @              $@      �?      @      �?      @                      �?      @              @      &@      @      @      @                      @      �?       @      �?      @      �?                      @              @rO  trP  bubhhubh)�rQ  }rR  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h<Kh=Kh>h"h#K �rS  h%�rT  RrU  (KK�rV  hV�C              �?rW  trX  bhJhZhEC       rY  �rZ  Rr[  h^Kh_h`Kh"h#K �r\  h%�r]  Rr^  (KK�r_  hE�C       r`  tra  bK�rb  Rrc  }rd  (hKhjMohkh"h#K �re  h%�rf  Rrg  (KMo�rh  hr�BHP         F                    �?0����?�           ��@                           �J@�-١�:�?]            @a@                          �>@     ��?,             P@������������������������       �                     �?                           �?�[|x��?+            �O@                          �T@r�q��?
             (@                          �P@����X�?             @������������������������       �                     @	       
                     E@�q�q�?             @������������������������       �                     �?                           @H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?�IєX�?!            �I@������������������������       �                     6@                          �W@ܷ��?��?             =@                           @I@�X�<ݺ?             2@                          �P@      �?              @                           �H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@                           �F@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @       =                     P@rr�J��?1            �R@       0                   �R@�G�z��?&             N@       #                    �?�q�q�?             B@       "                   �G@���}<S�?             7@        !                    �L@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     3@$       /                   �P@�θ�?
             *@%       .                    @O@r�q��?	             (@&       '                    �?z�G�z�?             $@������������������������       �                     @(       )                   �7@�q�q�?             @������������������������       �                      @*       +                    �K@      �?             @������������������������       �                     �?,       -                   �8@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?1       <                   �U@      �?             8@2       7                    @M@      �?             (@3       6                    �?�����H�?             "@4       5                    �K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @8       ;                   �U@�q�q�?             @9       :                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@>       E                   `V@؇���X�?             ,@?       D                   �L@$�q-�?
             *@@       A                    F@z�G�z�?             @������������������������       �                     @B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?G       �                    �?��Vu@z�?y           ��@H       o                    �G@X���o�?�            �u@I       Z                   @P@X~�pX��?.            @R@J       Y                   @K@PN��T'�?             ;@K       P                    �E@"pc�
�?             6@L       O                    �D@$�q-�?	             *@M       N                    @D@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @Q       R                    �F@�q�q�?             "@������������������������       �                     �?S       V                    @G@      �?              @T       U                    H@r�q��?             @������������������������       �                     �?������������������������       �                     @W       X                   @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @[       b                   @Q@��c:�?             G@\       a                    @F@�<ݚ�?             "@]       `                     E@�q�q�?             @^       _                     D@z�G�z�?             @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @c       h                   `U@4�B��?            �B@d       g                   �R@�����H�?             2@e       f                   `R@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     *@i       j                   @V@�\��N��?	             3@������������������������       �                      @k       n                    �D@��.k���?             1@l       m                    �B@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@������������������������       �                     @p       �                   @L@�`K?O��?�            `q@q       t                    @�����?r            �g@r       s                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     @u       �                   �I@HKS�l�?o            �f@v       �                     R@��)�G��?^            �c@w       �                    �O@XI�~�?\            @c@x       �                    �N@$�q-�?O            @`@y       �                   @C@�g+��@�?C            �[@z       �                   @@@���Ls�?'            @P@{       |                    6@�Ń��̧?             E@������������������������       �                     6@}       ~                    @L@P���Q�?             4@������������������������       �                     ,@       �                    �L@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �@@��<b���?             7@������������������������       �                     �?�       �                     L@"pc�
�?             6@�       �                   �B@�z�G��?             $@�       �                   �A@�<ݚ�?             "@������������������������       �                      @�       �                   @B@����X�?             @�       �                    �I@�q�q�?             @������������������������       �                      @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     �?�       �                   @B@�8��8��?             (@�       �                    �M@؇���X�?             @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     @�       �                   �F@��<b�ƥ?             G@�       �                   �E@���N8�?             5@������������������������       �        	             0@�       �                    �L@z�G�z�?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                     9@�       �                    .@�S����?             3@�       �                    @O@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    @O@@4և���?	             ,@������������������������       �                     @�       �                    E@ףp=
�?             $@������������������������       �                      @�       �                   @G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@�       �                    B@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @J@�+$�jP�?             ;@�       �                    �K@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                     O@�C��2(�?             6@������������������������       �                     &@�       �                   @K@"pc�
�?             &@�       �                     P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   �L@�VM�?5            @V@������������������������       �                     @�       �                    �L@�t����?4            @U@�       �                   �Y@nM`����?             G@�       �                    @J@��i#[�?             E@�       �                    @I@P���Q�?             4@�       �                    �H@�����H�?             "@������������������������       �                     @�       �                   `P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@�       �                    �K@�eP*L��?             6@�       �                    �J@      �?
             0@�       �                   �Q@      �?             @������������������������       �                     @������������������������       �                     @�       �                   �P@�z�G��?             $@�       �                   �O@؇���X�?             @������������������������       �                     @�       �                    @K@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    T@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @L@�q�q�?             @�       �                   �Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    U@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                     P@x�����?            �C@�       �                   `S@�r����?             >@�       �                    N@HP�s��?             9@�       �                   @M@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �M@���7�?             6@�       �                    @M@�����H�?             "@������������������������       �                      @�       �                   �O@؇���X�?             @������������������������       �                      @�       �                   �P@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     *@�       �                   �V@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   @P@X�<ݚ�?             "@������������������������       �                     @�       �                    `P@r�q��?             @�       �                   �R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�                          �?f���?�            �n@�                          @L@��s����?G            @Z@�                          �J@p`q�q��?5            �S@�                          @J@�^����?&            �M@�                         �W@�KM�]�?$            �L@�       �                    W@�S����?             C@�       �                    �B@l��\��?             A@�       �                     @@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    @F@XB���?             =@�       �                   `R@��S�ۿ?
             .@������������������������       �                     @�       �                    �E@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �        
             ,@                          �D@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@                        �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@                         @M@      �?             :@	                         �L@�z�G��?             $@
                        �P@      �?             @                         L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                        �S@�q�q�?             @                        �J@���Q��?             @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     �?                        �K@      �?
             0@������������������������       �                     @������������������������       �                     $@      0                  �I@B� ��?]            �a@      +                   @����>�?            �B@                        �;@¦	^_�?             ?@������������������������       �                     �?                         @G@������?             >@������������������������       �                      @                        �C@d}h���?             <@������������������������       �                      @      $                   @M@�z�G��?             4@       !                  @H@�����H�?             "@������������������������       �                     @"      #                  �H@      �?             @������������������������       �                     �?������������������������       �                     @%      &                   @N@�eP*L��?             &@������������������������       �                     @'      (                   �Q@      �?              @������������������������       �                     @)      *                   F@�q�q�?             @������������������������       �                      @������������������������       �                     �?,      -                  @G@r�q��?             @������������������������       �                     @.      /                   �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @1      f                   @����?C            �Y@2      M                   @L@�)V���?9            @V@3      4                   P@r�q��?&             N@������������������������       �                     ,@5      6                   �F@��<b���?             G@������������������������       �                     1@7      D                   @J@J�8���?             =@8      =                   T@X�<ݚ�?             2@9      <                   @G@      �?              @:      ;                  �R@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @>      C                   �I@z�G�z�?             $@?      @                  �X@�����H�?             "@������������������������       �                     @A      B                    H@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?E      F                   �J@"pc�
�?             &@������������������������       �                     @G      J                   @K@���Q��?             @H      I                  �T@�q�q�?             @������������������������       �                     �?������������������������       �                      @K      L                  �T@      �?              @������������������������       �                     �?������������������������       �                     �?N      ]                   @N@l��[B��?             =@O      T                  �S@�t����?             1@P      S                  �O@      �?              @Q      R                  �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @U      \                  �W@X�<ݚ�?             "@V      W                   T@�q�q�?             @������������������������       �                     �?X      Y                  �T@���Q��?             @������������������������       �                     �?Z      [                  �U@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     @^      _                  �R@      �?             (@������������������������       �                     @`      a                   �O@      �?              @������������������������       �                     �?b      c                   �P@և���X�?             @������������������������       �                     �?d      e                   S@�q�q�?             @������������������������       �                      @������������������������       �                     @g      l                   @O@����X�?
             ,@h      k                   @K@"pc�
�?             &@i      j                    I@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @m      n                    P@�q�q�?             @������������������������       �                      @������������������������       �                     �?ri  trj  bh�h"h#K �rk  h%�rl  Rrm  (KMoKK�rn  hV�B�        u@     �x@     �Y@     �A@      M@      @              �?      M@      @      $@       @      @       @      @              �?       @              �?      �?      �?      �?                      �?      @              H@      @      6@              :@      @      1@      �?      @      �?      �?      �?      �?                      �?      @              $@              "@       @      "@                       @     �F@      =@     �@@      ;@      (@      8@       @      5@       @       @               @       @                      3@      $@      @      $@       @       @       @      @              @       @       @               @       @              �?       @      �?              �?       @               @                      �?      5@      @      "@      @       @      �?      @      �?              �?      @              @              �?       @      �?      �?      �?                      �?              �?      (@              (@       @      (@      �?      @      �?      @              �?      �?      �?                      �?       @                      �?      m@     �v@     �Q@     �q@      7@      I@      @      7@      @      2@      �?      (@      �?      @              @      �?                      @      @      @      �?               @      @      �?      @      �?                      @      �?      �?              �?      �?                      @      3@      ;@      @       @      @       @      @      �?      @      �?      �?                      �?      @              (@      9@       @      0@       @      @              @       @                      *@      $@      "@       @               @      "@       @      "@       @                      "@      @             �G@     �l@      2@     `e@       @      @       @                      @      0@     �d@      &@      b@      $@      b@      $@      ^@      @      Z@      @     �M@      �?     �D@              6@      �?      3@              ,@      �?      @      �?                      @      @      2@      �?              @      2@      @      @       @      @               @       @      @       @      @               @       @       @              �?      �?              �?      &@      �?      @      �?       @              @              @      �?     �F@      �?      4@              0@      �?      @              @      �?      �?              9@      @      0@       @      @       @                      @      �?      *@              @      �?      "@               @      �?      �?      �?                      �?              8@      �?      �?              �?      �?              @      6@      @       @               @      @               @      4@              &@       @      "@       @      �?       @                      �?               @      =@      N@      @              9@      N@      1@      =@      *@      =@      �?      3@      �?       @              @      �?       @               @      �?                      &@      (@      $@      $@      @      @      @              @      @              @      @      @      �?      @              @      �?              �?      @              �?       @               @      �?               @      @      �?       @      �?                       @      �?       @               @      �?              @               @      ?@      @      :@       @      7@      �?       @               @      �?              �?      5@      �?       @               @      �?      @               @      �?      @      �?       @               @              *@       @      @       @                      @      @      @      @              �?      @      �?      �?      �?                      �?              @     `d@     �T@     @U@      4@      R@      @      J@      @     �I@      @      @@      @      ?@      @      @       @      @                       @      <@      �?      ,@      �?      @               @      �?       @                      �?      ,@              �?      @      �?                      @      3@              �?      �?              �?      �?              4@              *@      *@      @      @      �?      @      �?      �?              �?      �?                       @       @      @       @      @      �?      @      �?                      �?      $@      @              @      $@             �S@      O@      $@      ;@      "@      6@      �?               @      6@       @              @      6@               @      @      ,@      �?       @              @      �?      @      �?                      @      @      @      @               @      @              @       @      �?       @                      �?      �?      @              @      �?       @      �?                       @      Q@     �A@      P@      9@      I@      $@      ,@              B@      $@      1@              3@      $@      $@       @       @      @       @      �?              �?       @                      @       @       @       @      �?      @              @      �?      @                      �?              �?      "@       @      @              @       @       @      �?              �?       @              �?      �?              �?      �?              ,@      .@      @      (@      �?      @      �?       @               @      �?                      @      @      @      @       @      �?              @       @              �?      @      �?      �?               @      �?              @      "@      @      @              @      @      �?              @      @              �?      @       @               @      @              @      $@       @      "@       @      @              @       @                      @       @      �?       @                      �?ro  trp  bubhhubh)�rq  }rr  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h<Kh=Kh>h"h#K �rs  h%�rt  Rru  (KK�rv  hV�C              �?rw  trx  bhJhZhEC       ry  �rz  Rr{  h^Kh_h`Kh"h#K �r|  h%�r}  Rr~  (KK�r  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMMhkh"h#K �r�  h%�r�  Rr�  (KMM�r�  hr�B�H         �                    �?�+	G�?�           ��@                          �S@��4:���?�            Px@       J                   @L@ ˤ���?�            t@       5                   @G@�Cc}h��?�             l@       *                   �E@��cˣ��?a            �b@       )                   @C@|�9ǣ�?M            �]@                          @@@d۬����??            @W@                           �?@4և���?'             L@	       
                    5@r�q��?             @������������������������       �                     �?������������������������       �                     @                           @M@ "��u�?$             I@                           @L@ףp=
�?             >@������������������������       �                     3@                           &@���!pc�?             &@������������������������       �                     �?                           �L@z�G�z�?             $@                           :@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     4@                          �@@��G���?            �B@������������������������       �                     @       &                    `R@�t����?             A@                          �A@     ��?             @@������������������������       �                     "@                           @J@�LQ�1	�?             7@������������������������       �                      @       !                   @B@z�G�z�?
             .@                            �M@����X�?             @������������������������       �      �?             @������������������������       �                     @"       #                   �B@      �?              @������������������������       �                     �?$       %                    �K@؇���X�?             @������������������������       �                     �?������������������������       �                     @'       (                    B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     9@+       .                   @F@     ��?             @@,       -                    @M@      �?             @������������������������       �                      @������������������������       �      �?             @/       0       
             �?ȵHPS!�?             :@������������������������       �                     �?1       2                    @O@HP�s��?             9@������������������������       �                     5@3       4                    `P@      �?             @������������������������       �                      @������������������������       �                      @6       ;                    �?,N�_� �?6            �R@7       :                    J@؇���X�?             @8       9                    �P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @<       =                   �I@�L#���?/            �P@������������������������       �                     =@>       E                    �M@�KM�]�?             C@?       @                   �K@XB���?             =@������������������������       �                     2@A       B                    �G@�C��2(�?             &@������������������������       �                     "@C       D                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?F       I                    `P@�q�q�?             "@G       H                   �K@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @K       N                    �?R�L=��?:            @X@L       M                   �N@��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@O       t                    Q@fv�S��?2            �T@P       m                    @N@��U/��?#            �L@Q       Z                   @O@�L�lRT�?            �F@R       U                   �L@������?
             1@S       T                     M@�q�q�?             @������������������������       �                     �?������������������������       �                      @V       W                    �M@؇���X�?             ,@������������������������       �                     &@X       Y                   @M@�q�q�?             @������������������������       �                     �?������������������������       �                      @[       \                    P@և���X�?             <@������������������������       �                     �?]       l                    �M@�5��?             ;@^       i                   �P@      �?             6@_       b                   `P@�\��N��?             3@`       a                    �H@      �?              @������������������������       �                     �?������������������������       �                     �?c       h                    @K@��.k���?
             1@d       e                    @F@�q�q�?             (@������������������������       �                     @f       g                    �G@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @j       k                    �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @n       s                   @P@�8��8��?             (@o       p                    @P@z�G�z�?             @������������������������       �                      @q       r                   �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @u       v                   `R@HP�s��?             9@������������������������       �                      @w       ~                    �K@�t����?
             1@x       y                     G@�<ݚ�?             "@������������������������       �                     @z       {                    �J@�q�q�?             @������������������������       �                     �?|       }                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    X@�������?'             Q@�       �                    �?�Ƀ aA�?"            �M@�       �                   �V@*;L]n�?             >@�       �                    �O@�q�����?             9@�       �                    �E@���Q��?             4@������������������������       �                     @�       �                   `T@��.k���?             1@������������������������       �                     @�       �                    V@z�G�z�?             $@�       �                   �U@���Q��?             @�       �                    U@      �?             @�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   �U@�f7�z�?             =@�       �                    @J@�G��l��?             5@�       �                   �U@���!pc�?             &@������������������������       �                      @������������������������       �                     @�       �                     N@z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    �B@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?�����H�?             "@������������������������       �                     @�       �                    �D@r�q��?             @������������������������       �                     �?������������������������       �                     @�       
                   @L@bPD΂_�?�            �u@�       �                    �?��hJ,�?�            �m@�       �                    A@`<)�+�?-            @S@������������������������       �                     �?�       �                    �?P�Lt�<�?,             S@������������������������       �                     E@�       �                    S@�IєX�?             A@������������������������       �                     ,@�       �                   �U@ףp=
�?             4@������������������������       �                     �?�       �                   @X@�}�+r��?             3@�       �                    �H@ףp=
�?             $@�       �                    �F@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �                   `Q@���gb�?g             d@�       �                    @K@X�Cc�?#             L@�       �                   �D@p9W��S�?             C@�       �                    0@�q�q�?             @������������������������       �                     �?�       �                    =@z�G�z�?             @������������������������       �                     �?�       �                   @C@      �?             @�       �                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �H@     ��?             @@�       �                    @b�2�tk�?             2@�       �                    @G@     ��?
             0@�       �                   @P@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �        
             ,@�       �                   �P@      �?	             2@�       �                   @M@     ��?             0@�       �                    �?և���X�?             @������������������������       �                     �?�       �                   �K@�q�q�?             @�       �                    �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �N@�q�q�?             "@������������������������       �                      @�       �                   @O@և���X�?             @�       �                    @      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �E@(N:!���?D            @Z@�       �                   `Z@�nkK�?             G@�       �                    �?������?             B@�       �                    �B@�nkK�?             7@�       �                    �A@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �        	             ,@������������������������       �        	             *@�       �                   �Z@ףp=
�?             $@�       �                    �A@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       	                   @�:�B��?&            �M@�       �                    �?�k�'7��?%            �L@�       �                    �F@�J�4�?             9@�       �                   �W@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �J@�C��2(�?             6@������������������������       �                     *@�       �                   �[@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    �F@     ��?             @@������������������������       �                     @�       �                   @S@�<ݚ�?             ;@�       �                    @H@�q�q�?             @�       �                   �R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�                         `Z@r�q��?             8@�                         `T@�LQ�1	�?             7@�                           �H@      �?              @������������������������       �                     �?                         T@؇���X�?             @������������������������       �                     @������������������������       �                     �?                         @H@��S�ۿ?	             .@������������������������       �                      @                        �X@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         �?n�tl��?C            �Z@                         @z�G�z�?
             .@                         �N@�q�q�?             "@������������������������       �                     @                        �@@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @      &                  �I@�û��|�?9             W@                         @M@�חF�P�?             ?@������������������������       �                     @      %                   @�q�q�?             8@                         �?      �?             4@������������������������       �                      @                         �M@�E��ӭ�?             2@������������������������       �                      @                        �1@     ��?             0@                         �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         @C@$�q-�?	             *@������������������������       �                     @!      "                   �Q@؇���X�?             @������������������������       �                     @#      $                  �E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @'      F                   @Υf���?$            �N@(      ?                   U@�`���?            �H@)      :                   S@��J�fj�?            �B@*      1                   �?l��[B��?             =@+      .                   �L@�	j*D�?
             *@,      -                  �P@      �?             @������������������������       �                     �?������������������������       �                     @/      0                  @L@�����H�?             "@������������������������       �                     �?������������������������       �                      @2      3                   �N@     ��?	             0@������������������������       �                     @4      5                   @P@�eP*L��?             &@������������������������       �                      @6      7                    Q@�q�q�?             "@������������������������       �                     @8      9                   O@���Q��?             @������������������������       �                     @������������������������       �                      @;      <                   �M@      �?              @������������������������       �                     @=      >                  �S@      �?             @������������������������       �                     @������������������������       �                     �?@      A                   �?      �?             (@������������������������       �                     @B      C                   �L@�q�q�?             "@������������������������       �                      @D      E                   @N@؇���X�?             @������������������������       �                     @������������������������       �                     �?G      H                  �P@�q�q�?             (@������������������������       �                     @I      J                   @O@r�q��?             @������������������������       �                     @K      L                    P@�q�q�?             @������������������������       �                     �?������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMMKK�r�  hV�B�       `t@     �y@     �R@     �s@      E@     pq@      6@     @i@      1@     �`@      &@     �Z@      &@     �T@      @      J@      �?      @      �?                      @      @     �G@      @      ;@              3@      @       @      �?               @       @       @       @               @       @                      @              4@      @      >@      @              @      >@      @      =@              "@      @      4@               @      @      (@       @      @       @       @              @      �?      @              �?      �?      @      �?                      @      �?      �?              �?      �?                      9@      @      :@      @      @               @      @      �?      @      7@      �?               @      7@              5@       @       @       @                       @      @     @Q@      �?      @      �?       @               @      �?                      @      @     �O@              =@      @      A@      �?      <@              2@      �?      $@              "@      �?      �?      �?                      �?      @      @      @       @      @                       @              @      4@     @S@      �?      ,@      �?                      ,@      3@     �O@      1@      D@      0@      =@      @      *@       @      �?              �?       @               @      (@              &@       @      �?              �?       @              (@      0@      �?              &@      0@      &@      &@      $@      "@      �?      �?      �?                      �?      "@       @      @       @              @      @      @      @                      @      @              �?       @      �?                       @              @      �?      &@      �?      @               @      �?       @               @      �?                      @       @      7@               @       @      .@       @      @              @       @      �?      �?              �?      �?              �?      �?                       @     �@@     �A@      9@      A@      *@      1@      *@      (@       @      (@              @       @      "@              @       @       @      @       @      @      �?      �?      �?              �?      �?               @                      �?      @              @                      @      (@      1@      &@      $@      @       @               @      @               @       @       @                       @      �?      @      �?                      @       @      �?      @              @      �?              �?      @             `o@     �W@     `i@     �A@     �R@      @              �?     �R@       @      E@              @@       @      ,@              2@       @              �?      2@      �?      "@      �?      @      �?      @                      �?      @              "@              `@      @@      B@      4@      ;@      &@       @      @      �?              �?      @              �?      �?      @      �?       @               @      �?                      �?      9@      @      &@      @      &@      @      "@      �?      "@                      �?       @      @       @                      @               @      ,@              "@      "@      "@      @      @      @      �?               @      @       @      �?              �?       @                      @      @      @       @              @      @      @      @      @                      @      �?                       @     @W@      (@      F@       @     �A@      �?      6@      �?       @      �?       @                      �?      ,@              *@              "@      �?      �?      �?              �?      �?               @             �H@      $@     �G@      $@      5@      @      �?       @               @      �?              4@       @      *@              @       @      @                       @      :@      @      @              5@      @      �?       @      �?      �?              �?      �?                      �?      4@      @      4@      @      @       @              �?      @      �?      @                      �?      ,@      �?       @              @      �?      @                      �?              �?       @              H@     �M@      (@      @      @      @      @              @      @              @      @              @              B@      L@      @      :@              @      @      3@      @      .@               @      @      *@       @              @      *@       @      �?              �?       @              �?      (@              @      �?      @              @      �?      �?      �?                      �?              @      ?@      >@      8@      9@      5@      0@      ,@      .@      "@      @      �?      @      �?                      @       @      �?              �?       @              @      &@              @      @      @       @              @      @              @      @       @      @                       @      @      �?      @              @      �?      @                      �?      @      "@              @      @      @       @              �?      @              @      �?              @      @      @              �?      @              @      �?       @      �?                       @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMqhkh"h#K �r�  h%�r�  Rr�  (KMq�r�  hr�B�P         H                    �?6������?�           ��@       +                    �L@������?h            @d@                            �J@��#:���?G            �[@                           @D@�=C|F�?8            �U@       
                   �W@      �?
             0@       	                   �S@և���X�?             @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@                           �?h��@D��?.            �Q@                           @I@      �?             8@                           �G@�r����?             .@                           @G@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @                           �I@X�<ݚ�?             "@                           C@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @                           �?`Ql�R�?             �G@������������������������       �                     :@                           �G@���N8�?             5@                          `W@r�q��?             @������������������������       �                     @                            F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             .@!       $                    �?��+7��?             7@"       #                    U@      �?             @������������������������       �                     @������������������������       �                     �?%       &                    �?�S����?             3@������������������������       �                     *@'       *                   @M@      �?             @(       )                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @,       A                     P@��B����?!             J@-       4                   @O@�n_Y�K�?            �C@.       /                   �C@b�2�tk�?
             2@������������������������       �                     @0       3                    �?������?             .@1       2                   �G@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@5       >                    �?��s����?             5@6       =                    @O@      �?             0@7       8                    �N@ףp=
�?             $@������������������������       �                     @9       :                   `T@z�G�z�?             @������������������������       �                     @;       <                    U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @?       @                    �N@���Q��?             @������������������������       �                     @������������������������       �                      @B       G                    �P@$�q-�?             *@C       D                    `P@z�G�z�?             @������������������������       �                     �?E       F                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @I       �                   @M@���"�?x           ��@J       �                    �?V#L��?�            �p@K       L                    @���8�w�?�            @h@������������������������       �                     �?M       �                    �R@h2��v�?�             h@N       �                     P@��Y���?�            �g@O       P                   �:@�qE��E�?p            �d@������������������������       �                     ;@Q       �                    @O@�u����?`             a@R       s                   @F@�t`�4 �?V            �^@S       p                   �E@��� ��?*             O@T       o                   @C@lGts��?%            �K@U       \                   @@@��2(&�?             F@V       [                   �;@�IєX�?             1@W       X                    @L@r�q��?             @������������������������       �                     @Y       Z                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             &@]       ^                   �@@�+$�jP�?             ;@������������������������       �                      @_       `                    �E@H%u��?             9@������������������������       �                     �?a       n                    @L@�8��8��?             8@b       c                    @I@8�Z$���?	             *@������������������������       �                     @d       k                   �B@z�G�z�?             $@e       f                   �A@      �?              @������������������������       �                      @g       j                   @B@r�q��?             @h       i                    @K@      �?             @������������������������       �                      @������������������������       �      �?              @������������������������       �                      @l       m                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     &@q       r                    @M@����X�?             @������������������������       �                     @������������������������       ��q�q�?             @t       �                   @L@P���Q�?,             N@u       �                   �K@�1�`jg�?)            �K@v                            H@`Ӹ����?!            �F@w       |                   @I@      �?             0@x       {                    H@ףp=
�?             $@y       z                    @F@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @}       ~                    @G@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     =@�       �                    �G@ףp=
�?             $@������������������������       �                      @�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �?@������?
             .@������������������������       �                     �?�       �                   �I@d}h���?	             ,@�       �                    F@8�Z$���?             *@������������������������       �                     @�       �                   @G@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@�       �                    B@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     E@:PZ(8?�?1            @R@������������������������       �                     @�       �                    @K@(���X�?/            @Q@�       �                    �J@8�A�0��?             6@�       �                    �?�����?             3@�       �                    �I@r�q��?             @������������������������       �                     @�       �                    A@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @G@$�q-�?             *@�       �                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     @�       �                    @��|�5��?             �G@�       �                    �?�������?             F@�       �                    <@@4և���?             ,@�       �                   �:@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                   �I@������?             >@�       �                   �G@��<b���?             7@�       �                    C@�q�q�?             .@�       �                    �P@      �?              @�       �                    �N@z�G�z�?             @������������������������       �                      @�       �                    $@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �E@և���X�?             @������������������������       �                     �?�       �                   �F@      �?             @������������������������       �                     �?�       �                    �N@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   �K@և���X�?             @�       �                     P@      �?             @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �H@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       X                   �M@�.7,]�?�            s@�                          �?NB�!��?�            @o@�                         @[@���|���?8             V@�       �                    @J@8�$�>�?6            �U@�       �                   `X@�rF���?!            �K@�       �                   @W@ \� ���?            �H@�       �                   �R@z�G�z�?             D@�       �                    �F@�d�����?             3@������������������������       �                     (@�       �                   @P@����X�?             @������������������������       �                     �?�       �                   `Q@�q�q�?             @�       �                    �G@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                   �U@�����?             5@������������������������       �                     &@�       �                    �G@z�G�z�?             $@�       �                    �D@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �B@X�<ݚ�?             "@������������������������       �                      @�       �                   �W@և���X�?             @������������������������       �                     �?�       �                    @E@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �J@�P�*�?             ?@�       �                    P@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @K@X�<ݚ�?             ;@�       �                   �O@�q�q�?             @������������������������       �                     �?�       �                   @T@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �K@�ՙ/�?             5@������������������������       �                      @�       �                    �L@D�n�3�?             3@�       �                    @L@      �?              @�       �                   �Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    U@���Q��?             @������������������������       �                     �?�       �                   @Y@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @M@�eP*L��?             &@������������������������       �                     �?�       �                   �O@���Q��?             $@������������������������       �                      @                         �U@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                      @      K                   @�����?h            @d@      H                  �\@�ӖF2��?^            �a@      /                   @L@��L��d�?\            @a@                         �E@��ϭ�*�?M             ]@                         @B@�(\����?             D@	                         �?@4և���?             ,@
                         �A@�C��2(�?	             &@������������������������       �                      @                         X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     :@                         @S@h�˹�?2             S@                        �P@z�G�z�?             >@������������������������       �        
             .@                         �?���Q��?	             .@                         �H@�z�G��?             $@                         R@���Q��?             @������������������������       �                     @������������������������       �                      @                         R@z�G�z�?             @                         Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         �F@���Q��?             @������������������������       �                      @������������������������       �                     @!      *                   Y@���.�6�?             G@"      )                   @I@�?�|�?            �B@#      (                   W@�IєX�?             1@$      %                   �?      �?             @������������������������       �                     �?&      '                   @H@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     *@������������������������       �                     4@+      .                   �I@�<ݚ�?             "@,      -                  �Y@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @0      G                   Y@8�A�0��?             6@1      B                   V@�ՙ/�?             5@2      A                   @M@��S���?
             .@3      >                  �T@��
ц��?	             *@4      9                   �?X�<ݚ�?             "@5      8                   �L@z�G�z�?             @6      7                  �P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @:      ;                   �L@      �?             @������������������������       �                     �?<      =                  @R@�q�q�?             @������������������������       �                      @������������������������       �                     �??      @                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @C      D                   �?r�q��?             @������������������������       �                     �?E      F                  �W@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     �?I      J                  `]@      �?             @������������������������       �                     @������������������������       �                     �?L      W                  @Z@      �?
             4@M      N                   �D@X�Cc�?             ,@������������������������       �                      @O      R                  �P@      �?             (@P      Q                  @O@      �?             @������������������������       �                      @������������������������       �                      @S      T                  �U@      �?              @������������������������       �                     @U      V                   �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @Y      \                   �?�2�o�U�?             �K@Z      [                  �N@`2U0*��?             9@������������������������       �                     �?������������������������       �                     8@]      ^                   �?��S���?             >@������������������������       �                     @_      d                   �N@� �	��?             9@`      c                   @      �?              @a      b                  @P@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?e      j                   �O@j���� �?	             1@f      g                   @      �?             @������������������������       �                     �?h      i                  �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @k      p                  �T@��
ц��?             *@l      o                   @�<ݚ�?             "@m      n                   S@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMqKK�r�  hV�B       �t@     �x@      ^@      E@     @W@      1@      S@      &@      (@      @      @      @      @      �?              �?      @                      @      "@              P@      @      2@      @      *@       @      @       @      @                       @      @              @      @      @      @      @                      @       @              G@      �?      :@              4@      �?      @      �?      @              �?      �?      �?                      �?      .@              1@      @      �?      @              @      �?              0@      @      *@              @      @      �?      @              @      �?               @              ;@      9@      .@      8@      &@      @              @      &@      @       @      @       @                      @      "@              @      1@      �?      .@      �?      "@              @      �?      @              @      �?      �?      �?                      �?              @      @       @      @                       @      (@      �?      @      �?      �?              @      �?              �?      @               @             �j@     Pv@     �D@     @l@      1@      f@      �?              0@      f@      .@      f@      .@     �b@              ;@      .@     �^@      &@     �[@       @      K@      @     �H@      @      C@      �?      0@      �?      @              @      �?       @      �?                       @              &@      @      6@       @              @      6@      �?               @      6@       @      &@              @       @       @      �?      @               @      �?      @      �?      @               @      �?      �?               @      �?      �?      �?                      �?              &@              &@       @      @              @       @      �?      @     �L@      @      J@       @     �E@       @      ,@      �?      "@      �?      @              @      �?                      @      �?      @              @      �?                      =@      �?      "@               @      �?      �?      �?                      �?              @      @      &@      �?              @      &@       @      &@              @       @      @       @                      @      �?                      ;@      �?      �?              �?      �?              8@     �H@      @              4@     �H@      "@      *@      @      *@      @      �?      @              �?      �?              �?      �?              �?      (@      �?      @      �?                      @              "@      @              &@      B@      "@     �A@      �?      *@      �?      �?              �?      �?                      (@       @      6@      @      2@      @      $@      �?      @      �?      @               @      �?       @               @      �?                      @      @      @      �?              @      @              �?      @       @      @                       @               @      @      @      @      �?      �?      �?      �?                      �?       @                      @       @      �?              �?       @             �e@     ``@     �c@     @W@      @@      L@      >@      L@      (@     �E@      (@     �B@      @     �@@      @      ,@              (@      @       @      �?              @       @      @       @      @                       @      �?               @      3@              &@       @       @       @       @               @       @                      @      @      @       @              @      @              �?      @      @              @      @                      @      2@      *@      @      �?              �?      @              .@      (@       @      @      �?              �?      @              @      �?              *@       @       @              &@       @      @      @       @      �?       @                      �?      @       @              �?      @      �?      @                      �?      @      @              �?      @      @               @      @       @      @                       @       @             @_@     �B@      ^@      6@     �]@      3@     �Z@      $@     �C@      �?      *@      �?      $@      �?       @               @      �?              �?       @              @              :@             �P@      "@      8@      @      .@              "@      @      @      @      @       @      @                       @      @      �?      �?      �?      �?                      �?      @               @      @       @                      @     �E@      @      B@      �?      0@      �?      @      �?      �?               @      �?      �?              �?      �?      *@              4@              @       @       @       @               @       @              @              *@      "@      *@       @       @      @      @      @      @      @      @      �?       @      �?       @                      �?       @              �?      @              �?      �?       @               @      �?              �?      @              @      �?               @              @      �?      �?              @      �?       @      �?       @                      �?      �?      @              @      �?              @      .@      @      "@       @              @      "@       @       @               @       @              �?      @              @      �?       @      �?                       @              @      1@      C@      �?      8@      �?                      8@      0@      ,@      @              &@      ,@      �?      @      �?      @      �?                      @              �?      $@      @      @      �?      �?               @      �?              �?       @              @      @      @       @       @       @               @       @              @                      @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJQY%hG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMChkh"h#K �r�  h%�r�  Rr�  (KMC�r�  hr�B�F         B       	             �?�Z���?�           ��@       %                    �?      �?d             e@       "                    U@      �?&            �Q@                           5@�f7�z�?!             M@������������������������       �                      @                          �A@��>4և�?              L@������������������������       �                     @       !                    �P@
j*D>�?             J@	                           �J@`�(c�?            �H@
                            E@\X��t�?             7@������������������������       �                     @                           �H@�����?             3@������������������������       �                     @                           �I@և���X�?             ,@                           @I@���Q��?             $@������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     @                           S@�θ�?             :@                          �G@�IєX�?             1@                           �O@      �?             @                          @F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     *@                            �O@X�<ݚ�?             "@                          `T@z�G�z�?             @������������������������       �                     @                           �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @#       $                   �V@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?&       '                    @H@@4և���?>            �X@������������������������       �                     =@(       1                    @I@�θV�?,            @Q@)       0                   �T@���|���?             &@*       +                   �O@�q�q�?             @������������������������       �                     �?,       -                    �H@z�G�z�?             @������������������������       �                      @.       /                    Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @2       5                    C@�8���?%             M@3       4                     @      �?              @������������������������       �                     �?������������������������       �                     �?6       A                   �Q@h�����?#             L@7       8                    �N@HP�s��?             9@������������������������       �        	             *@9       :                    �?r�q��?             (@������������������������       �                     @;       <                   @F@�<ݚ�?             "@������������������������       �                     @=       >                    �O@�q�q�?             @������������������������       �                     �??       @                     Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ?@C       �                    �?�=`��?w           ��@D       �                   @L@d4(x���?�            �t@E       v                   @C@|)���?�            @j@F       s                    `R@H%u��?A             Y@G       r                     P@��l��??            @X@H       M                     I@�=C|F�?9            �U@I       J                   @B@�IєX�?             1@������������������������       �                     *@K       L                    �E@      �?             @������������������������       �                     �?������������������������       �                     @N       Q                    @؇���X�?2            �Q@O       P                     @      �?              @������������������������       �                     �?������������������������       �                     �?R       S                    +@�G�V�e�?0             Q@������������������������       �                      @T       W                    �J@R���Q�?)             N@U       V                   @@@և���X�?             @������������������������       �                     @������������������������       �                     @X       Y                    .@���C��?$            �J@������������������������       �                      @Z       q                   @B@�:�]��?#            �I@[       j                   �A@�����?             E@\       ]                    5@      �?             @@������������������������       �                      @^       c                    8@�8��8��?             8@_       `                     L@�q�q�?             @������������������������       �                     �?a       b                    @N@      �?              @������������������������       �                     �?������������������������       �                     �?d       e                   �=@���N8�?             5@������������������������       �                     @f       i                   �?@@4և���?             ,@g       h                    �O@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @k       l                    @K@z�G�z�?             $@������������������������       �                      @m       n                    @L@      �?              @������������������������       �      �?              @o       p                    �M@r�q��?             @������������������������       �z�G�z�?             @������������������������       �                     �?������������������������       �                     "@������������������������       �                     $@t       u                    B@�q�q�?             @������������������������       �                      @������������������������       �                     �?w       �                    �H@���7�?I            �[@x       �                    @H@ףp=
�?             >@y       �                   �J@ 	��p�?             =@z                           J@      �?             0@{       |                    @G@��S�ۿ?             .@������������������������       �        	             &@}       ~                   @I@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?�       �                    @L@�(\����?4             T@������������������������       �                    �@@�       �                   �I@`�q�0ܴ?            �G@������������������������       �                    �@@�       �                   @J@؇���X�?
             ,@������������������������       �                      @������������������������       �                     (@�       �                   �R@P&��?O            �]@�       �                    �H@F�����?&            �L@�       �                   �O@�E��ӭ�?             2@������������������������       �                      @�       �                    @F@     ��?	             0@�       �                   @Q@���Q��?             @�       �                     E@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                    �M@�q�q�?            �C@�       �                    @M@
j*D>�?             :@�       �                   �P@��Q��?             4@�       �                    �J@������?
             .@������������������������       �                      @�       �                   @M@և���X�?             @������������������������       �                     �?�       �                    �L@�q�q�?             @�       �                    @K@z�G�z�?             @�       �                   �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    Q@���Q��?             @������������������������       �                      @�       �                    @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �P@�q�q�?             @�       �                   �M@z�G�z�?             @������������������������       �                      @�       �                   �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                     P@8�Z$���?	             *@������������������������       �                      @�       �                    `P@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �Z@�jTM��?)            �N@�       �                   �S@����>4�?'             L@�       �                   �R@��S�ۿ?             .@������������������������       �                     �?�       �                   `S@@4և���?             ,@�       �                    �J@$�q-�?
             *@������������������������       �                      @�       �                    �K@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �D@���?            �D@������������������������       �                     (@�       �                     G@J�8���?             =@������������������������       �                     @�       �                   `T@�+e�X�?             9@������������������������       �                     @�       �                   �W@�����?             5@�       �                    @K@�r����?             .@������������������������       �                     @�       �                     N@      �?              @�       �                     M@�q�q�?             @������������������������       �                     �?�       �                   �U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                     M@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?ҳ�wY;�?�            �m@�       �                    @L@�C+����?@            @Y@�       �                    ;@$��$�L�?3            �S@������������������������       �                     �?�       �                   @\@�:�^���?2            �S@�       �                    �B@�S(��d�?1            @S@�       �                   �V@�	j*D�?	             *@�       �                   �T@z�G�z�?             @�       �                   `R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   `Q@      �?(             P@�       �                    @K@�C��2(�?             6@������������������������       �                     0@�       �                   �P@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     E@������������������������       �                     �?�       �                    Q@���|���?             6@�       �                   @L@؇���X�?	             ,@������������������������       �                      @�       �                    �M@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   @T@      �?              @������������������������       �                     @�       �                    @M@      �?             @������������������������       �                      @������������������������       �                      @�                         �N@���<��?^             a@�                          @����S��?%             M@�       �                    @G@J��D��?"             K@������������������������       �                     @�       
                   �N@t�F�}�?            �I@�       �                   �?@�MI8d�?            �B@�       �                    @M@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �F@؇���X�?            �A@������������������������       �                      @�                          @K@�+$�jP�?             ;@�                            I@      �?              @������������������������       �                     @������������������������       �                     @                        �G@�KM�]�?             3@������������������������       �                     �?                         J@�X�<ݺ?
             2@������������������������       �                     *@      	                  �K@z�G�z�?             @                         �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        �F@և���X�?	             ,@                          R@�q�q�?             "@                        �9@      �?              @                         $@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         P@ܩ�d	��?9            �S@������������������������       �                      @                         @E@����O��?3            �Q@                         @      �?             0@������������������������       �        
             ,@                         �B@      �?              @������������������������       �                     �?������������������������       �                     �?      *                   �I@���|���?'            �K@      %                    H@�\��N��?             3@                          �E@���!pc�?             &@������������������������       �                     �?!      "                   �F@z�G�z�?             $@������������������������       �                     @#      $                   T@����X�?             @������������������������       �                      @������������������������       �                     @&      '                  �S@      �?              @������������������������       �                     @(      )                   @I@      �?             @������������������������       �                     @������������������������       �                     �?+      B                    Q@�E��ӭ�?             B@,      ?                  `X@��R[s�?            �A@-      >                    O@�n`���?             ?@.      3                  @S@��+7��?             7@/      0                   �J@      �?             @������������������������       �                     �?1      2                  �P@���Q��?             @������������������������       �                      @������������������������       �                     @4      5                   T@@�0�!��?             1@������������������������       �                     @6      7                  `U@      �?	             (@������������������������       �                      @8      9                  �U@ףp=
�?             $@������������������������       �                     @:      =                  `V@r�q��?             @;      <                   �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @@      A                   �L@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMCKK�r�  hV�B0        u@     �x@     �_@      E@     �A@     �A@      8@      A@       @              6@      A@              @      6@      >@      3@      >@      *@      $@              @      *@      @      @               @      @      @      @      @       @              @      @              @      4@      �?      0@      �?      @      �?      �?              �?      �?                       @              *@      @      @      �?      @              @      �?      �?              �?      �?              @              @              &@      �?      &@                      �?     �V@      @      =@              O@      @      @      @       @      @      �?              �?      @               @      �?       @               @      �?              @             �K@      @      �?      �?              �?      �?              K@       @      7@       @      *@              $@       @      @              @       @      @              �?       @              �?      �?      �?      �?                      �?      ?@             �j@      v@      M@     �p@      1@      h@      (@      V@      &@     �U@      &@      S@      �?      0@              *@      �?      @      �?                      @      $@      N@      �?      �?              �?      �?              "@     �M@               @      "@     �I@      @      @              @      @              @     �G@       @              @     �G@      @      C@       @      >@               @       @      6@      �?       @              �?      �?      �?      �?                      �?      �?      4@              @      �?      *@      �?      @              @      �?                      @       @       @               @       @      @      �?      �?      �?      @      �?      @              �?              "@              $@      �?       @               @      �?              @     @Z@      @      ;@       @      ;@       @      ,@      �?      ,@              &@      �?      @              @      �?              �?                      *@      �?               @     �S@             �@@       @     �F@             �@@       @      (@       @                      (@     �D@     @S@      :@      ?@      *@      @               @      *@      @       @      @       @      �?       @                      �?               @      &@              *@      :@      &@      .@      @      *@      @      &@               @      @      @              �?      @       @      @      �?       @      �?       @                      �?       @                      �?      @       @       @              �?       @      �?                       @      @       @      @      �?       @               @      �?              �?       @                      �?       @      &@               @       @      @       @                      @      .@      G@      &@     �F@      �?      ,@              �?      �?      *@      �?      (@               @      �?      @      �?                      @              �?      $@      ?@              (@      $@      3@      @              @      3@      @               @      3@       @      *@              @       @      @       @      �?      �?              �?      �?      �?                      �?              @              @      @      �?              �?      @             @c@      U@     �S@      6@     �Q@       @              �?     �Q@      @     �Q@      @      "@      @      �?      @      �?      �?              �?      �?                      @       @              O@       @      4@       @      0@              @       @      @                       @      E@                      �?       @      ,@       @      (@               @       @      @              @       @              @       @      @               @       @               @       @             �R@      O@      1@     �D@      1@     �B@      @              ,@     �B@      @      ?@      �?      �?              �?      �?              @      >@               @      @      6@      @      @              @      @               @      1@      �?              �?      1@              *@      �?      @      �?      �?      �?                      �?              @       @      @      @      @       @      @       @      �?              �?       @                      @      �?              @                      @      M@      5@       @              I@      5@      .@      �?      ,@              �?      �?              �?      �?             �A@      4@      "@      $@       @      @              �?       @       @      @              @       @               @      @              �?      @              @      �?      @              @      �?              :@      $@      :@      "@      9@      @      1@      @      @      @      �?               @      @       @                      @      ,@      @      @              "@      @               @      "@      �?      @              @      �?      �?      �?      �?                      �?      @               @              �?      @      �?                      @              �?r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ��fbhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMihkh"h#K �r�  h%�r�  Rr�  (KMi�r�  hr�B�N         �                    �?�#i����?�           ��@       !       	             �?D�X%��?           �x@                            `P@X�<ݚ�?$             K@                          �T@���Q��?"             I@       
                    �H@r٣����?            �@@                           �D@X�<ݚ�?             "@������������������������       �                     @       	                   �F@r�q��?             @������������������������       �                     �?������������������������       �                     @                           �N@      �?             8@                            N@@�0�!��?             1@                           ;@@4և���?	             ,@������������������������       �                     �?������������������������       �                     *@                          �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                          �V@�t����?             1@                           @M@�θ�?             *@������������������������       �                      @                           �N@���Q��?             @������������������������       �                     �?                           U@      �?             @������������������������       �                     �?                          �U@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �X@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @"       W                    @I@yF�?�            �u@#       2                    �D@Nṧ'
�?>            �W@$       %                   �O@�����H�?             ;@������������������������       �                     "@&       )                    �B@r�q��?             2@'       (                   �U@�q�q�?             @������������������������       �                      @������������������������       �                     �?*       +                    @C@�r����?             .@������������������������       �                     @,       /                    �C@z�G�z�?	             $@-       .                   �Q@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?0       1                   @Q@؇���X�?             @������������������������       �                     �?������������������������       �                     @3       F                    �G@ҳ�wY;�?)             Q@4       E                    @G@X�<ݚ�?             B@5       @                   �T@      �?             @@6       ;                    H@�㙢�c�?             7@7       8                    @F@���!pc�?             &@������������������������       �                     @9       :                   @E@���Q��?             @������������������������       �                      @������������������������       �                     @<       =                    �F@�8��8��?
             (@������������������������       �                     @>       ?                   @O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?A       B                    �E@�����H�?             "@������������������������       �                     @C       D                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @G       P                    �H@      �?             @@H       O                   `Y@z�G�z�?
             .@I       J                    @H@$�q-�?	             *@������������������������       �                     @K       L                    J@؇���X�?             @������������������������       �                     @M       N                   �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @Q       R                   �L@�t����?             1@������������������������       �                     "@S       V                   �Q@      �?              @T       U                   �O@r�q��?             @������������������������       �                      @������������������������       �      �?             @������������������������       �                      @X       �                    `P@T���RB�?�             o@Y       �                    �O@ ��(��?�            @l@Z       �                   @M@����B"�?�             i@[       n                   �<@ ����?X            @`@\       i                   �9@z�G�z�?             9@]       ^                     L@�KM�]�?             3@������������������������       �                     @_       f                    5@؇���X�?             ,@`       a                    �N@�8��8��?	             (@������������������������       �                     @b       e                    @O@r�q��?             @c       d                    '@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @g       h                   �7@      �?              @������������������������       �                     �?������������������������       �                     �?j       k                     L@      �?             @������������������������       �                      @l       m                    �L@      �?             @������������������������       �                      @������������������������       �      �?              @o       �                   �I@�#-���?E            @Z@p                          @F@p��@���?5            @U@q       |                   �E@�q��/��?             G@r       u                    �I@��p\�?            �D@s       t                   �?@      �?              @������������������������       �                     �?������������������������       �                     �?v       {                    �K@�7��?            �C@w       x                    @K@8�Z$���?             *@������������������������       �                      @y       z                   @B@���Q��?             @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     :@}       ~                    @M@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @�       �                    @O@ ���J��?            �C@������������������������       �                    �B@�       �                   @G@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @L@R���Q�?             4@������������������������       �                     $@�       �                   �J@�z�G��?             $@������������������������       �                      @�       �                    @M@      �?              @������������������������       �                     @�       �                    �M@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �K@�ګH9�?)            �Q@�       �                   @P@և���X�?             <@������������������������       �                      @�       �                    @J@�n_Y�K�?             :@������������������������       �                      @�       �                    @K@X�<ݚ�?             2@�       �                   �Q@�eP*L��?             &@�       �                   �P@؇���X�?             @������������������������       �                     @�       �                   �P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �R@����X�?             @�       �                   �Q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    N@(L���?            �E@������������������������       �                     �?�       �                    R@���H��?             E@������������������������       �        
             ,@�       �                    �M@�>4և��?             <@�       �                   �U@     ��?             0@�       �                   `T@���Q��?             $@�       �                    @L@      �?              @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                      @�       �                   �Y@r�q��?             @������������������������       �                     @�       �                     M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@�       �                     P@`�Q��?             9@�       �                    ;@������?	             .@������������������������       �                     @�       �                   �?@���|���?             &@������������������������       �                      @�       �                   �I@�<ݚ�?             "@������������������������       �                     @�       �                   �K@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �M@���Q��?             $@������������������������       �                     @�       �                   �R@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     7@�                          �K@,Tg�x0�?�             u@�       �                   @C@T�6|���?             j@�       �                    �?����X�?             @�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     F@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �T@pLBQh��?y             i@�       �                    �?r�q��?<             X@�       �                    �?��hJ,�?             A@������������������������       �                     .@�       �                   �R@�d�����?	             3@�       �                   `P@��S�ۿ?             .@������������������������       �                     @�       �                    @G@      �?              @������������������������       �                     @�       �                    @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @�n`���?'             O@�       �                    Q@���5��?$            �L@�       �                    �H@ ��WV�?             :@�       �                   �K@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@�       �                   �Q@�n`���?             ?@������������������������       �                     �?�       �                    �?r�q��?             >@������������������������       �        
             0@�       �                    �J@X�Cc�?	             ,@�       �                    @G@�����H�?             "@������������������������       �                     @�       �                     I@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @K@z�G�z�?             @�       �                   @S@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�                          @����?=            @Z@�       �                    �?b �57�?;            �Y@�       �                   �W@������?             B@������������������������       �        
             2@�       �                    �?�X�<ݺ?
             2@������������������������       �                     @�       �                    �F@$�q-�?             *@������������������������       �                     "@�       �                    @I@      �?             @������������������������       �                     �?������������������������       �                     @�                          �?�qM�R��?'            �P@�                          �G@�����H�?             B@�                          �U@`2U0*��?             9@�       �                    @@@�q�q�?             @������������������������       �                     �?�       �                    @C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@                         W@���!pc�?             &@������������������������       �                     @                         �H@և���X�?             @                         Y@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @	      
                  `Z@`Jj��?             ?@������������������������       �                     9@                          G@�q�q�?             @������������������������       �                     @������������������������       �                      @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?      <                  @M@     ^�?Q             `@            
             �?�q�q�?"            �I@                         �Q@�n_Y�K�?             *@                        @C@      �?              @                         �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @                         �R@���Q��?             @������������������������       �                     @������������������������       �                      @      %                    N@�I�w�"�?             C@                        �G@X�<ݚ�?             "@������������������������       �                      @      $                   @����X�?             @       !                  �I@�q�q�?             @������������������������       �                     @"      #                   �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?&      1                    P@д>��C�?             =@'      (                   �?��S�ۿ?	             .@������������������������       �                     @)      *                   �N@ףp=
�?             $@������������������������       �                     @+      0                   @O@؇���X�?             @,      /                  �=@      �?             @-      .                   $@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @2      ;                   @R@����X�?
             ,@3      :                   @      �?              @4      5                   �P@և���X�?             @������������������������       �                     �?6      7                  �C@      �?             @������������������������       �                      @8      9                    Q@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @=      B      	             �?���!pc�?/            @S@>      A                  @R@P���Q�?             4@?      @                   P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             2@C      F                  �P@���dQ'�?$            �L@D      E                   �M@      �?
             0@������������������������       �                      @������������������������       �                     ,@G      L                  `Q@�>$�*��?            �D@H      I                   Q@؇���X�?             @������������������������       �                     @J      K                   �?      �?             @������������������������       �                     �?������������������������       �                     @M      N                   �L@ҳ�wY;�?             A@������������������������       �                      @O      ^                   �N@��
ц��?             :@P      ]                   @��S���?             .@Q      \                   �M@��
ц��?	             *@R      Y                   @M@�q�q�?             (@S      V                   �?X�<ݚ�?             "@T      U                  @T@      �?             @������������������������       �                     @������������������������       �                     �?W      X                   V@���Q��?             @������������������������       �                      @������������������������       �                     @Z      [                   W@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @_      d                   S@���|���?             &@`      c                   @���Q��?             @a      b                  �R@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?e      h                   �P@r�q��?             @f      g                  @U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMiKK�r�  hV�B�       `u@     �x@     �V@     0s@      8@      >@      4@      >@       @      9@      @      @              @      @      �?              �?      @              @      5@      @      ,@      �?      *@      �?                      *@       @      �?       @                      �?              @      (@      @      $@      @       @               @      @              �?       @       @      �?              �?       @               @      �?               @       @               @       @              @             �P@     Pq@      ;@      Q@      @      8@              "@      @      .@      �?       @               @      �?               @      *@              @       @       @      �?       @      �?      �?              �?      �?      @      �?                      @      8@      F@      0@      4@      (@      4@      @      3@      @       @              @      @       @               @      @              �?      &@              @      �?      @              @      �?               @      �?      @              �?      �?      �?                      �?      @               @      8@      @      (@      �?      (@              @      �?      @              @      �?       @      �?                       @       @              @      (@              "@      @      @      @      �?       @              @      �?               @      D@      j@      D@     @g@      @@      e@      ,@      ]@      @      4@       @      1@              @       @      (@      �?      &@              @      �?      @      �?      �?              �?      �?                      @      �?      �?      �?                      �?      @      @               @      @      �?       @              �?      �?      "@      X@      @     �S@      @     �D@      @      C@      �?      �?              �?      �?               @     �B@       @      &@               @       @      @       @       @              �?              :@       @      @               @       @      �?      �?      C@             �B@      �?      �?      �?                      �?      @      1@              $@      @      @       @              �?      @              @      �?      @      �?                      @      2@     �J@      (@      0@       @              $@      0@               @      $@       @      @      @      �?      @              @      �?       @      �?                       @      @              @       @       @       @       @                       @      @              @     �B@      �?              @     �B@              ,@      @      7@      @      &@      @      @       @      @               @       @      @       @              �?      @              @      �?       @               @      �?                      (@       @      1@      @      &@              @      @      @       @               @      @              @       @       @       @                       @      @      @              @      @      �?      @                      �?              7@     `o@     @U@     @f@      >@       @      @      �?      �?              �?      �?              �?      @      �?                      @      f@      9@     �S@      1@      =@      @      .@              ,@      @      ,@      �?      @              @      �?      @              �?      �?              �?      �?                      @      I@      (@      I@      @      9@      �?      @      �?              �?      @              2@              9@      @              �?      9@      @      0@              "@      @       @      �?      @              @      �?              �?      @              �?      @      �?       @               @      �?                       @              @     @X@       @      X@      @     �A@      �?      2@              1@      �?      @              (@      �?      "@              @      �?              �?      @             �N@      @      @@      @      8@      �?       @      �?      �?              �?      �?              �?      �?              6@               @      @      @              @      @      �?      @              @      �?              @              =@       @      9@              @       @      @                       @      �?      �?      �?                      �?     @R@     �K@      1@      A@       @      @      @       @       @       @               @       @              @               @      @              @       @              "@      =@      @      @       @               @      @       @      @              @       @      �?       @                      �?              �?      @      8@      �?      ,@              @      �?      "@              @      �?      @      �?      @      �?      �?              �?      �?                       @              @      @      $@      @      @      @      @      �?              @      @               @      @      �?              �?      @                      �?              @      L@      5@      3@      �?      �?      �?      �?                      �?      2@             �B@      4@      ,@       @               @      ,@              7@      2@      �?      @              @      �?      @      �?                      @      6@      (@       @              ,@      (@      @       @      @      @      @      @      @      @      @      �?      @                      �?       @      @       @                      @       @      �?       @                      �?              �?               @      @      @       @      @      �?      @      �?                      @      �?              @      �?      �?      �?              �?      �?              @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ$�phG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r   tr  bK�r  Rr  }r  (hKhjMWhkh"h#K �r  h%�r  Rr  (KMW�r  hr�BK         :                    �?"��G,�?�           ��@       +                    �?� ��fd�?a            @b@       
                    C@�eP*L��?$            �K@                           8@���!pc�?             &@������������������������       �                     @                          �@@      �?              @������������������������       �                      @       	                    �H@r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @                           �H@�zv�X�?             F@                           X@���|���?             &@                           T@X�<ݚ�?             "@                          �P@����X�?             @                            F@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                           �C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @       *                     Q@:ɨ��?            �@@       #                   `T@r֛w���?             ?@                          �G@�LQ�1	�?             7@                          �E@      �?              @������������������������       �                     �?������������������������       �                     �?       "                    �J@�����?             5@       !                    R@�q�q�?             @                            �I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     .@$       %                    @M@      �?              @������������������������       �                     @&       '                    �N@���Q��?             @������������������������       �                      @(       )                   �V@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @,       3                    �N@x��B�R�?=            �V@-       2                   �P@ ��ʻ��?/             Q@.       /                   `P@      �?             0@������������������������       �                     *@0       1                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        $             J@4       5                    @@���}<S�?             7@������������������������       �                     �?6       9                   @R@���7�?             6@7       8                    @O@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                     &@;       �                    �I@V��f_�?]           `�@<       =                    �@@�Z����?v            `h@������������������������       �                     &@>       I                    �B@��*(��?o             g@?       B                    �?ҳ�wY;�?             1@@       A                    @B@      �?             @������������������������       �                     @������������������������       �                     �?C       H                    @�θ�?
             *@D       G                    V@r�q��?	             (@E       F                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?J       w                    �?�:�>��?b            �d@K       R                    �D@��0%�?4            �V@L       Q                    �C@�8��8��?             8@M       P                   @T@      �?              @N       O                    @C@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     0@S       v                   �Y@.��<�?)            �P@T       q                    �H@r�q��?&             N@U       n                    @H@     ��?             H@V       i                   �V@�T|n�q�?            �E@W       X                    @F@������?            �B@������������������������       �                     (@Y       Z                   @E@�J�4�?             9@������������������������       �                     "@[       \                    H@      �?             0@������������������������       �                     �?]       h                   �R@z�G�z�?             .@^       g                   `R@      �?	             (@_       f                   @Q@"pc�
�?             &@`       a                    @G@      �?              @������������������������       �                     @b       e                    �G@�q�q�?             @c       d                   @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @j       k                    �E@      �?             @������������������������       �                      @l       m                   �X@      �?             @������������������������       �                     �?������������������������       �                     @o       p                    J@���Q��?             @������������������������       �                     @������������������������       �                      @r       s                   �M@�8��8��?             (@������������������������       �                     @t       u                    S@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @x       y                   �E@�d�����?.             S@������������������������       �                     "@z       �                    �?�iޤ��?)            �P@{       �                    �G@ףp=
�?             >@|       }                    �E@P���Q�?             4@������������������������       �                     "@~       �                    @F@�C��2(�?             &@       �                   �U@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @H@z�G�z�?             $@�       �                   �V@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �F@��%��?            �B@�       �                   �Z@8�Z$���?             *@������������������������       �                     $@�       �                    @C@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �G@      �?             8@�       �                   �Y@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                   �I@��S���?	             .@������������������������       �                      @�       �                    @��
ц��?             *@�       �                   �S@      �?             (@������������������������       �                     @�       �                    @H@�q�q�?             "@������������������������       �                     @�       �                    �H@      �?             @������������������������       �                      @�       �                    U@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     �?�                          �M@~y���?�            �x@�       �                    �?v����?            @i@�       �                    R@"pc�
�?P            �`@�       �                    @Ԫ2��?A            �\@������������������������       �                      @�       �                   �A@      �?@             \@������������������������       �                     @@�       �                   @C@z�G�z�?0             T@�       �                    �J@X�Cc�?             ,@������������������������       �                      @�       �                   @B@�q�q�?             (@�       �                    @K@�z�G��?             $@������������������������       �                     �?�       �                    @L@�<ݚ�?             "@������������������������       �                     @������������������������       ����Q��?             @������������������������       �                      @�       �                    @L@�U�=���?)            �P@�       �                    @K@���7�?             F@�       �                    �J@�>����?             ;@������������������������       �        	             *@�       �                    L@؇���X�?	             ,@������������������������       �                     $@�       �                    P@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     1@�       �                    �L@��2(&�?             6@�       �                   @K@      �?              @�       �                   @H@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     ,@�       �                    @J@X�<ݚ�?             2@������������������������       �                     @�       �                   �R@��S���?             .@������������������������       �                      @�       �                   �S@��
ц��?             *@�       �                    �K@z�G�z�?             @�       �                    @K@�q�q�?             @������������������������       �                     �?�       �                   �R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �U@      �?              @������������������������       �                     @�       �                   �Y@���Q��?             @������������������������       �                      @�       �                     M@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @L@��
P��?/            �Q@�       �                   �T@֭��F?�?            �G@�       �                    �?X�<ݚ�?             B@�       �                   �8@؇���X�?             ,@������������������������       �                     �?�       �                    Q@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?�       �                    @���|���?             6@�       �                    �J@�z�G��?             4@������������������������       �                     @�       �                    �K@ҳ�wY;�?
             1@�       �                   `Q@���Q��?             $@�       �                    @K@z�G�z�?             @������������������������       �                     �?�       �                   @M@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �I@����X�?             @������������������������       �                     @�       �                   �N@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    @"pc�
�?	             &@�       �                    @K@�<ݚ�?             "@�       �                    �?�q�q�?             @�       �                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @J@      �?             @�       �                   @Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�                          @8����?             7@�                          @M@�q�q�?             5@�                          �?������?             1@�                           �L@����X�?             @�       �                   �P@      �?             @������������������������       �                     �?������������������������       �                     @                         H@�q�q�?             @������������������������       �                      @������������������������       �                     �?                         �L@z�G�z�?             $@                         V@      �?              @������������������������       �                     �?������������������������       �                     �?      	                  @R@      �?              @������������������������       �                     @
                        `U@      �?              @������������������������       �                     �?������������������������       �                     �?                        @D@      �?             @������������������������       �                      @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @      *                   �N@�P��Af�?h            �g@      !                   �?؇���X�?            �H@                        @E@ףp=
�?             >@������������������������       �        	             *@                          @N@@�0�!��?
             1@                         K@���!pc�?             &@                         H@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?                        @O@      �?              @                        �L@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @"      )                  �P@���y4F�?
             3@#      &                   @N@���|���?             &@$      %                  @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?'      (                   F@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @+      8                   �?����?K            �a@,      7                  �?@Ћ����?,            �T@-      4                  �=@�S����?
             3@.      3                   @O@      �?             0@/      2                   4@z�G�z�?             @0      1                   '@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     &@5      6                   �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        "            �O@9      V                   �R@��S���?             N@:      M                   @6C�z��?            �L@;      B                  @J@��c:�?             G@<      A                  �E@�C��2(�?             6@=      >                   �?      �?              @������������������������       �                     �??      @                  �C@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     ,@C      D                   �O@�q�q�?             8@������������������������       �                     $@E      F                   �?      �?             ,@������������������������       �                     @G      L                    Q@�z�G��?             $@H      I                   �P@      �?             @������������������������       �                     �?J      K                   S@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @N      O                   �O@"pc�
�?             &@������������������������       �                     �?P      Q                    P@ףp=
�?             $@������������������������       �                     @R      U                   �P@؇���X�?             @S      T                   T@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @r	  tr
  bh�h"h#K �r  h%�r  Rr  (KMWKK�r  hV�Bp       @s@     �z@     @\@     �@@      9@      >@       @      @      @              @      @               @      @      �?      @               @      �?      1@      ;@      @      @      @      @      @       @      @      �?              �?      @              �?      �?              �?      �?                       @       @              $@      7@       @      7@      @      4@      �?      �?              �?      �?               @      3@       @      @       @      �?              �?       @                      @              .@      @      @      @               @      @               @       @      �?       @                      �?       @              V@      @     �P@      �?      .@      �?      *@               @      �?       @                      �?      J@              5@       @              �?      5@      �?      $@      �?              �?      $@              &@             `h@     �x@     @X@     �X@      &@             �U@     �X@      &@      @      �?      @              @      �?              $@      @      $@       @      @       @               @      @              @                      �?     �R@      W@      3@      R@       @      6@       @      @       @      @               @       @      �?              @              0@      1@      I@      $@      I@      "@     �C@      @      B@      @     �@@              (@      @      5@              "@      @      (@      �?              @      (@      @      "@       @      "@       @      @              @       @      �?      �?      �?              �?      �?              �?                      @      �?                      @      @      @       @              �?      @      �?                      @       @      @              @       @              �?      &@              @      �?      @      �?                      @      @              L@      4@      "@             �G@      4@      ;@      @      3@      �?      "@              $@      �?      @      �?              �?      @              @               @       @      @       @      @                       @      @              4@      1@      &@       @      $@              �?       @               @      �?              "@      .@      �?       @               @      �?               @      @       @              @      @      @      @              @      @      @      @              @      @               @      @      �?      �?               @      �?              �?     �X@     pr@      N@     �a@      8@      [@      0@     �X@       @              ,@     �X@              @@      ,@     �P@      "@      @       @              @      @      @      @              �?      @       @      @              @       @               @      @     �N@       @      E@       @      9@              *@       @      (@              $@       @       @       @                       @              1@      @      3@      @      @      @      �?              �?      @                      @              ,@       @      $@              @       @      @       @              @      @      �?      @      �?       @              �?      �?      �?              �?      �?                       @      @      @      @               @      @               @       @      �?              �?       @              B@      A@      =@      2@      4@      0@      (@       @              �?      (@      �?      (@                      �?       @      ,@      @      ,@              @      @      &@      @      @      @      �?      �?              @      �?              �?      @                      @       @      @              @       @       @       @                       @       @              "@       @      @       @      @       @      �?      �?      �?                      �?      @      �?      �?      �?      �?                      �?       @              @               @              @      0@      @      ,@      @      *@       @      @      �?      @      �?                      @      �?       @               @      �?               @       @      �?      �?              �?      �?              �?      @              @      �?      �?      �?                      �?      @      �?       @              �?      �?      �?                      �?               @      C@      c@      @      E@      @      ;@              *@      @      ,@      @       @       @      �?      �?      �?      �?              �?      @      �?      @              @      �?                      @              @      @      .@      @      @      �?       @               @      �?              @      @              @      @                       @      ?@     �[@      @     �S@      @      0@      �?      .@      �?      @      �?      �?              �?      �?                      @              &@       @      �?              �?       @                     �O@      <@      @@      <@      =@      3@      ;@       @      4@       @      @              �?       @      @              @       @                      ,@      1@      @      $@              @      @      @              @      @      @      @              �?      @       @               @      @                      @      "@       @              �?      "@      �?      @              @      �?      @      �?      @                      �?      @                      @r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJW:+LhG        hNhG        h<Kh=Kh>h"h#K �r  h%�r  Rr  (KK�r  hV�C              �?r  tr  bhJhZhEC       r  �r  Rr  h^Kh_h`Kh"h#K �r  h%�r  Rr  (KK�r  hE�C       r   tr!  bK�r"  Rr#  }r$  (hKhjMehkh"h#K �r%  h%�r&  Rr'  (KMe�r(  hr�BN         �                   @M@�#i����?�           ��@       ]                    �?p�L���?�            `s@                           -@H0sE�d�?�             l@       	                    *@���N8�?             5@                           �M@�C��2(�?	             &@                           @L@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @
                           @O@���Q��?             $@                           �N@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           �?@��Y��?�            �i@                          �G@z�G�z�?             4@                            M@X�<ݚ�?             "@                           8@����X�?             @������������������������       �                     �?                          �C@r�q��?             @                           @H@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                      @������������������������       �                     &@       6                    @L@̫��+�?~             g@                           �E@`Ӹ����?;            �V@������������������������       �        
             0@       -                   @J@@-�_ .�?1            �R@                            @J@Pa�	�?+            �P@������������������������       �                     @@!       $                    �J@�IєX�?             A@"       #                    E@      �?              @������������������������       �                     �?������������������������       �                     �?%       &                   �A@      �?             @@������������������������       �        	             1@'       ,                    �K@��S�ۿ?             .@(       )                    @K@�����H�?             "@������������������������       �                     @*       +                    F@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �                     @.       /                   �J@      �?              @������������������������       �                     �?0       1                   �K@؇���X�?             @������������������������       �                      @2       3                    �G@z�G�z�?             @������������������������       �                      @4       5                   �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @7       P                   �I@$�3c�s�?C            �W@8       A                    @M@�L���?5            �R@9       >                    �L@z�G�z�?             .@:       =                   �>@ףp=
�?             $@;       <                    5@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @?       @                   �?@���Q��?             @������������������������       ��q�q�?             @������������������������       �                      @B       G                   @@@����˵�?*            �M@C       D                   �>@؇���X�?
             ,@������������������������       �                     &@E       F                    @O@�q�q�?             @������������������������       �                     �?������������������������       �                      @H       O                    @N@����?�?             �F@I       J                    �M@@4և���?
             ,@������������������������       �                     "@K       L                    D@z�G�z�?             @������������������������       �                     �?M       N                   �G@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     ?@Q       \                    @P@      �?             4@R       S                   �J@X�Cc�?
             ,@������������������������       �                      @T       W                   �K@      �?             (@U       V                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?X       Y                    @M@z�G�z�?             $@������������������������       �                     @Z       [                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @^       i                    �?k�q��?7            @U@_       h                    `Q@�c�Α�?             =@`       g                    C@�<ݚ�?             ;@a       f                    :@�eP*L��?             &@b       e                   �8@      �?              @c       d                   �7@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �        
             0@������������������������       �                      @j       s                    �?��X��?'             L@k       p                   �>@ҳ�wY;�?
             1@l       o                    �M@r�q��?             @m       n                   �8@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @q       r                    @O@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?t       �                   �J@:�&���?            �C@u       v                   �D@��a�n`�?             ?@������������������������       �                     "@w       z                   �E@��2(&�?             6@x       y                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?{       |                   @H@�}�+r��?             3@������������������������       �                     "@}       �                   �H@ףp=
�?             $@~                           �J@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                     Q@      �?              @�       �                    �K@z�G�z�?             @������������������������       �                      @�       �                     O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       "                   �L@������?
           �z@�       �                    �?z�G��?�             t@�       �                    �?P�;�&��?8            @U@�       �                    �A@��}*_��?             ;@������������������������       �                      @�       �                    @I@`�Q��?             9@�       �                   �V@�8��8��?             (@������������������������       �                     "@�       �                    X@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @L@��
ц��?             *@�       �                    �J@�z�G��?             $@�       �                    �I@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �? 	��p�?(             M@������������������������       �                    �A@�       �                    @�㙢�c�?             7@�       �                   �T@��s����?             5@�       �                    @I@X�<ݚ�?             "@�       �                    �H@�q�q�?             @�       �                   �R@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        
             (@������������������������       �                      @�                          @J@(���@��?�            `m@�       �                    @H@�JX-��?k            @f@�       �                    �?x�=���?S            �a@�       �                   �W@v ��?            �E@�       �                    �F@���|���?            �@@�       �                    �C@��+7��?             7@�       �                    @C@      �?             $@������������������������       �                     @�       �                   �Q@����X�?             @������������������������       �r�q��?             @������������������������       �                     �?�       �                     E@$�q-�?             *@������������������������       �                     @�       �                    �E@؇���X�?             @�       �                    S@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �R@���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                   �Y@z�G�z�?             $@�       �                    �D@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   @P@z�09JX�?9            @X@������������������������       �                     ,@�       �                   `T@�?a/��?3            �T@�       �                   @S@և���X�?             5@�       �                    �?�q�q�?             2@�       �                   �P@���Q��?             $@������������������������       �                      @�       �                    �E@      �?              @������������������������       �                     @�       �                    R@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �F@      �?              @������������������������       �                     @�       �                   �R@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    Y@���-T��?&             O@�       �                    @B@`Jj��?             ?@�       �                    �?����X�?             @�       �                    �A@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     8@�       �                   �Y@��a�n`�?             ?@�       �                    �G@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    @H%u��?             9@������������������������       �                     4@�       �                   @Z@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �V@�\��N��?             C@�       �                    �?��H�}�?             9@�       �                   �R@X�<ݚ�?             2@�       �                    @I@���|���?             &@�       �                   `P@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?r�q��?             @�       �                    O@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    @I@؇���X�?             @������������������������       �                     @�       �                   �S@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?�	j*D�?             *@������������������������       �                     �?�       �                    @I@      �?             (@�       �                   �X@���Q��?             @������������������������       �                     @������������������������       �                      @�                          @Y@؇���X�?             @������������������������       �                     @������������������������       �                     �?                         �J@P̏����?#            �L@                         �?؇���X�?             @                        �P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                         @L@�-���?             I@	                        �T@      �?             D@
                        �P@�q�q�?             >@                         @K@8�Z$���?	             *@                         �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @                         �K@��.k���?	             1@                         @K@     ��?             0@                         �?      �?             @������������������������       �                     �?������������������������       �                     @                        �R@      �?             (@������������������������       �                     @                         �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@      !                   Z@�z�G��?             $@                         �Q@      �?              @                        �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @#      `                    P@��
ц��?D             Z@$      =                   �?���Q��?<            �V@%      <                  �Y@���V��?             �F@&      /      	             �?��2(&�?             F@'      (                   �N@r�q��?             2@������������������������       �                     @)      .                  `T@      �?	             (@*      +                  �R@ףp=
�?             $@������������������������       �                     @,      -                   �O@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @0      ;                  �V@ȵHPS!�?             :@1      :                   �M@��2(&�?             6@2      9                  `S@      �?              @3      4                   @M@����X�?             @������������������������       �                      @5      6                  �O@���Q��?             @������������������������       �                      @7      8                  �P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             ,@������������������������       �                     @������������������������       �                     �?>      ?                   �?�L�lRT�?            �F@������������������������       �                      @@      A                  @N@��J�fj�?            �B@������������������������       �                      @B      I                  �Q@���Q��?            �A@C      H                   �N@ףp=
�?             $@D      E                   �M@r�q��?             @������������������������       �                      @F      G                  �P@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @J      [                   @�q�����?             9@K      P                   �?D�n�3�?             3@L      O                   V@      �?             @M      N                   @M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @Q      Z                   �O@��S���?	             .@R      W                   V@�n_Y�K�?             *@S      V                  �T@�<ݚ�?             "@T      U                   T@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @X      Y                   @M@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                      @\      _                  �T@r�q��?             @]      ^                   S@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @a      d                   S@؇���X�?             ,@b      c                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@r)  tr*  bh�h"h#K �r+  h%�r,  Rr-  (KMeKK�r.  hV�BP       `u@     �x@     �O@     �n@      8@      i@      @      0@      �?      $@      �?      @              @      �?                      @      @      @      @      �?              �?      @                      @      3@      g@      @      0@      @      @       @      @      �?              �?      @      �?      @              �?      �?       @               @       @                      &@      .@      e@      @     �U@              0@      @     �Q@       @      P@              @@       @      @@      �?      �?      �?                      �?      �?      ?@              1@      �?      ,@      �?       @              @      �?      @      �?       @               @              @       @      @      �?              �?      @               @      �?      @               @      �?       @      �?                       @      &@     �T@      @      Q@      @      (@      �?      "@      �?      @              @      �?                      @       @      @       @      �?               @      @      L@       @      (@              &@       @      �?              �?       @              �?      F@      �?      *@              "@      �?      @              �?      �?      @      �?       @              �?              ?@      @      .@      @      "@       @              @      "@      �?      �?              �?      �?               @       @              @       @      @       @                      @              @     �C@      G@      5@       @      5@      @      @      @      @      @       @      @       @                      @      @                      @      0@                       @      2@      C@      &@      @      �?      @      �?      �?              �?      �?                      @      $@      �?      $@                      �?      @      @@      @      <@              "@      @      3@       @      �?       @                      �?      �?      2@              "@      �?      "@      �?      @      �?                      @              @      @      @      �?      @               @      �?       @      �?                       @      @             pq@      b@     �l@     @V@     �Q@      ,@      1@      $@               @      1@       @      &@      �?      "@               @      �?              �?       @              @      @      @      @      @      @              @      @                      @      @              K@      @     �A@              3@      @      1@      @      @      @       @      @       @      �?       @                      �?              @      @              (@               @              d@     �R@     @]@     �N@     �X@     �D@      4@      7@      (@      5@      @      1@      @      @              @      @       @      @      �?              �?      �?      (@              @      �?      @      �?       @               @      �?                      @      @      @      @                      @       @       @      @       @               @      @              @             �S@      2@      ,@             @P@      2@      (@      "@      (@      @      @      @               @      @       @      @              �?       @      �?                       @      @       @      @               @       @               @       @                      @     �J@      "@      =@       @      @       @      @       @      @                       @      �?              8@              8@      @       @      @              @       @              6@      @      4@               @      @       @                      @      2@      4@      "@      0@       @      $@      @      @       @      @              @       @              @      �?      @      �?              �?      @               @              �?      @              @      �?              �?      @              @      �?       @               @      �?              "@      @              �?      "@      @      @       @      @                       @      @      �?      @                      �?     �E@      ,@      @      �?       @      �?              �?       @              @             �B@      *@      >@      $@      4@      $@      &@       @      @       @               @      @               @              "@       @      "@      @      @      �?              �?      @              @      @              @      @       @      @                       @              �?      $@              @      @      @      �?      �?      �?      �?                      �?      @                       @      H@      L@      B@      K@      @      C@      @      C@      @      .@              @      @      "@      �?      "@              @      �?      @              @      �?               @              @      7@      @      3@      @      @       @      @               @       @      @               @       @      �?       @                      �?      �?                      ,@              @      �?              =@      0@       @              5@      0@               @      5@      ,@      "@      �?      @      �?       @              @      �?      @                      �?      @              (@      *@      &@       @      @      �?      �?      �?              �?      �?               @               @      @       @      @      @       @       @       @       @                       @      @              �?      @      �?       @              �?               @      �?      @      �?       @               @      �?                      @      (@       @      �?       @               @      �?              &@        r/  tr0  bubhhubh)�r1  }r2  (hhh	h
hNhKhKhG        hh hNhJF<KdhG        hNhG        h<Kh=Kh>h"h#K �r3  h%�r4  Rr5  (KK�r6  hV�C              �?r7  tr8  bhJhZhEC       r9  �r:  Rr;  h^Kh_h`Kh"h#K �r<  h%�r=  Rr>  (KK�r?  hE�C       r@  trA  bK�rB  RrC  }rD  (hKhjM]hkh"h#K �rE  h%�rF  RrG  (KM]�rH  hr�BXL         J                    �?�#i����?�           ��@       )                    �L@�zœ���?e            `c@                           �G@n����W�?C            �X@                          @W@�ʈD��?            �E@       
                   �V@8�Z$���?             :@       	                    @D@�8��8��?             8@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     2@������������������������       �                      @������������������������       �                     1@       (                    �K@d}h���?(             L@                          �A@ \� ���?$            �H@                           9@r�q��?             @������������������������       �                     �?������������������������       �                     @       '                   �T@�T|n�q�?             �E@       "                    �I@     ��?             @@                           �?�q�q�?             2@                           O@և���X�?             @                           �H@z�G�z�?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                      @       !                   �S@���!pc�?             &@                           �?�����H�?             "@������������������������       �                     @                           �H@z�G�z�?             @������������������������       �                     @                            @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @#       &                   �N@@4և���?
             ,@$       %                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     &@������������������������       �                     @*       G                    `P@��>4և�?"             L@+       0                    @M@�Q����?             D@,       /                    T@�q�q�?             @-       .                    P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @1       <                    �?�ʻ����?             A@2       3                    @N@���N8�?             5@������������������������       �                     @4       5                   �E@X�Cc�?	             ,@������������������������       �                      @6       9                    �O@�q�q�?             (@7       8                   @M@      �?              @������������������������       �                      @������������������������       �                     @:       ;                   �R@      �?             @������������������������       �                     �?������������������������       �                     @=       F                   @R@�θ�?	             *@>       ?                    �N@      �?             @������������������������       �                     �?@       E                    P@���Q��?             @A       D                    @�q�q�?             @B       C                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @H       I                   `V@      �?
             0@������������������������       �        	             .@������������������������       �                     �?K       �                    �?�^��[i�?k           �@L       y                   �I@h������?�            �r@M       N                   �:@`Jj��?g            `c@������������������������       �                     ?@O       p                    @N@6uH���?Q             _@P       g                   @F@���W���?8            �U@Q       Z                    @L@�㙢�c�?              G@R       U                    �E@�>����?             ;@S       T                    @D@�q�q�?             @������������������������       �                      @������������������������       �                     �?V       W                   �A@ �q�q�?             8@������������������������       �                     &@X       Y                    @K@$�q-�?	             *@������������������������       �                     &@������������������������       �      �?              @[       d                    �M@�����?             3@\       c                   @B@����X�?
             ,@]       ^                    �L@���Q��?             $@������������������������       �                     �?_       b                   �@@�q�q�?             "@`       a                    =@z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @������������������������       �      �?             @������������������������       �                     @e       f                    D@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @h       o                   @G@�(\����?             D@i       j                   �F@�}�+r��?             3@������������������������       �                     @k       n                    �H@      �?
             0@l       m                    @F@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                     5@q       x                   �?@P�Lt�<�?             C@r       s                    �O@r�q��?             @������������������������       �                     �?t       w                    �P@z�G�z�?             @u       v                   �=@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @@z       �                    @E@����6Z�?_            `b@{       |                    @D@`2U0*��?             9@������������������������       �        
             (@}       �                    �D@$�q-�?             *@~                          �P@�C��2(�?             &@������������������������       �                     @�       �                    S@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �P@<�yr��?N            �^@�       �                    @N@���Q��?+            @P@�       �                    �E@�`���?            �H@������������������������       �                     @�       �                    �H@��S���?            �F@������������������������       �                     @�       �                   @L@��
ц��?            �C@�       �                    @L@r�q��?             (@������������������������       �                     "@�       �                    K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    P@�5��?             ;@�       �                   @M@      �?             (@�       �                    �M@      �?             @������������������������       �                      @������������������������       �                      @�       �                   @O@      �?              @�       �                   @N@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   `P@��S���?             .@������������������������       �                     �?�       �                    �K@      �?             ,@�       �                     J@r�q��?             @������������������������       ��q�q�?             @������������������������       �                     @�       �                    �M@      �?              @������������������������       �                     @������������������������       �                      @�       �                   �N@      �?             0@������������������������       �                     "@�       �                     P@����X�?             @������������������������       �                     @�       �                   @P@�q�q�?             @������������������������       �                     �?�       �                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �S@�MWl��?#            �L@�       �                   �R@HP�s��?             9@�       �                    �K@8�Z$���?	             *@�       �                    R@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `R@�C��2(�?             &@������������������������       �                     "@�       �                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                   `T@     ��?             @@������������������������       �                     @�       �                   @[@�<ݚ�?             ;@�       �                   �W@���B���?             :@�       �                   �V@������?
             .@�       �                    @L@8�Z$���?	             *@�       �                    �J@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@������������������������       �                      @�       �                    �G@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?�                          @N@�W��?�            Pq@�       �                   �:@��X��?4             U@�       �                    �N@      �?             0@������������������������       �                     $@�       �                     Q@r�q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    $@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �E@h+�v:�?,             Q@�       �                    @X�<ݚ�?             2@�       �                    �?      �?             0@�       �                    A@�q�q�?             "@������������������������       �                     @�       �                   �C@      �?             @�       �                     L@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     �?�       �                     P@և���X�?             @������������������������       �                     @�       �                    D@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �F@`�Q��?              I@������������������������       �                      @�       �                     K@�q�q�?             H@�       �                     I@      �?             ,@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �I@�������?             A@�       �                    �?�㙢�c�?             7@������������������������       �                      @�       �                   �G@������?             .@�       �                    �Q@�q�q�?             @�       �                     P@z�G�z�?             @�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                   �J@�eP*L��?             &@������������������������       �                      @�       �                     Q@�q�q�?             "@�       �                    �?      �?              @�       �                   �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �K@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                         �E@Pu�����?q             h@                         @C@�.ߴ#�?"            �N@                         �A@ �Cc}�?             <@                         R@���7�?             6@������������������������       �                     �?������������������������       �                     5@                         W@�q�q�?             @������������������������       �                     �?	      
                  �Z@z�G�z�?             @������������������������       �                     @                         @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �@@                         P@�X����?O            �`@                         @K@���7�?             6@������������������������       �                     *@                          M@�����H�?             "@                         @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @      ,                   �?bOvj6��?C            �[@      +                   V@"pc�
�?            �@@                        �Q@����X�?             5@                        �P@؇���X�?             @                        �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @      &                  �S@X�Cc�?	             ,@       #                  `R@X�<ݚ�?             "@!      "                    K@      �?              @������������������������       �                     �?������������������������       �                     �?$      %                   �H@և���X�?             @������������������������       �                     @������������������������       �                     @'      (                   U@z�G�z�?             @������������������������       �                     �?)      *                   �J@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             (@-      T                   @�eP*L��?+            @S@.      9                   S@Pa�.l�?&            �P@/      0                   �F@�t����?             1@������������������������       �                      @1      2                    J@z�G�z�?
             .@������������������������       �                     @3      4                   �J@���!pc�?             &@������������������������       �                     �?5      6                   �M@z�G�z�?             $@������������������������       �                     @7      8                  @Q@�q�q�?             @������������������������       �                      @������������������������       �                     @:      =                   �G@�w��#��?             I@;      <                  �V@�q�q�?             @������������������������       �                     @������������������������       �                      @>      S                   �P@v�X��?             F@?      @                   T@�q�q�?            �C@������������������������       �                     "@A      B                  �T@*;L]n�?             >@������������������������       �                     @C      R                  �Y@$��m��?             :@D      O                  `W@�q�q�?             8@E      F                  �T@���Q��?	             .@������������������������       �                     @G      H                  @U@      �?             (@������������������������       �                     @I      J                   �I@�q�q�?             "@������������������������       �                      @K      L                   V@؇���X�?             @������������������������       �                     @M      N                    L@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @P      Q                    M@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @U      \                  �W@���Q��?             $@V      W                   S@      �?              @������������������������       �                     �?X      Y                   �L@և���X�?             @������������������������       �                      @Z      [                   �N@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @rI  trJ  bh�h"h#K �rK  h%�rL  RrM  (KM]KK�rN  hV�B�       `u@     �x@     @]@      C@     �T@      0@     �C@      @      6@      @      6@       @      @       @               @      @              2@                       @      1@              F@      (@     �B@      (@      �?      @      �?                      @      B@      @      9@      @      (@      @      @      @      @      �?      @              �?      �?               @       @      @       @      �?      @              @      �?      @              �?      �?              �?      �?                       @      *@      �?       @      �?              �?       @              &@              &@              @              A@      6@      3@      5@      @       @      �?       @      �?                       @      @              .@      3@      @      0@              @      @      "@               @      @      @       @      @       @                      @      @      �?              �?      @              $@      @      @      @      �?               @      @       @      �?      �?      �?              �?      �?              �?                       @      @              .@      �?      .@                      �?      l@      v@      I@     �o@      $@      b@              ?@      $@     �\@      "@     @S@       @      C@       @      9@      �?       @               @      �?              �?      7@              &@      �?      (@              &@      �?      �?      @      *@      @      $@      @      @      �?              @      @      �?      @      �?       @               @       @       @              @       @      @               @       @      �?      �?     �C@      �?      2@              @      �?      .@      �?      @              @      �?                      &@              5@      �?     �B@      �?      @              �?      �?      @      �?      @              @      �?                      �?              @@      D@     �Z@      �?      8@              (@      �?      (@      �?      $@              @      �?      @      �?                      @               @     �C@     �T@      :@     �C@      8@      9@              @      8@      5@      @              2@      5@       @      $@              "@       @      �?       @                      �?      0@      &@      "@      @       @       @       @                       @      @      �?      @      �?      @                      �?      @              @       @              �?      @      @      �?      @      �?       @              @      @       @      @                       @       @      ,@              "@       @      @              @       @      �?      �?              �?      �?      �?                      �?      *@      F@       @      7@       @      &@      �?      �?              �?      �?              �?      $@              "@      �?      �?      �?                      �?              (@      &@      5@      @              @      5@      @      5@      @      &@       @      &@       @       @               @       @                      "@       @              �?      $@      �?                      $@      �?             �e@     �Y@      ;@     �L@      �?      .@              $@      �?      @      �?       @              �?      �?      �?              �?      �?                      @      :@      E@      $@       @      $@      @      @      @      @              @      @       @      @      �?              �?      @      �?              @      @      @              �?      @              @      �?                       @      0@      A@               @      0@      @@      @      @      �?      @      �?                      @      @              "@      9@      @      3@               @      @      &@      @       @      @      �?      �?      �?      �?                      �?      @                      �?              "@      @      @       @              @      @       @      @      �?       @               @      �?              �?      @      �?                      @      �?             �b@     �F@      M@      @      9@      @      5@      �?              �?      5@              @       @              �?      @      �?      @              �?      �?      �?                      �?     �@@             �V@      E@      5@      �?      *@               @      �?      �?      �?      �?                      �?      @             @Q@     �D@      ;@      @      .@      @      @      �?      �?      �?      �?                      �?      @              "@      @      @      @      �?      �?      �?                      �?      @      @              @      @              @      �?      �?              @      �?      @                      �?      (@              E@     �A@      C@      =@      @      (@       @              @      (@              @      @       @      �?               @       @              @       @      @       @                      @     �@@      1@       @      @              @       @              ?@      *@      :@      *@      "@              1@      *@              @      1@      "@      1@      @      "@      @      @              @      @              @      @      @               @      @      �?      @               @      �?      �?              �?      �?       @      �?       @                      �?               @      @              @      @      @      @              �?      @      @       @               @      @              @       @                       @rO  trP  bubhhubh)�rQ  }rR  (hhh	h
hNhKhKhG        hh hNhJؽ�hG        hNhG        h<Kh=Kh>h"h#K �rS  h%�rT  RrU  (KK�rV  hV�C              �?rW  trX  bhJhZhEC       rY  �rZ  Rr[  h^Kh_h`Kh"h#K �r\  h%�r]  Rr^  (KK�r_  hE�C       r`  tra  bK�rb  Rrc  }rd  (hKhjMChkh"h#K �re  h%�rf  Rrg  (KMC�rh  hr�B�F         �                    �?�/�$�y�?�           ��@       '       	             �?@�0�!��?�            px@                           �J@      �?&             P@                          �T@�P�*�?             ?@                            E@�eP*L��?             6@������������������������       �                     @       
                   �G@      �?             0@       	                   �>@؇���X�?             @������������������������       �                     �?������������������������       �                     @                           Q@X�<ݚ�?             "@                           �H@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          �V@�����H�?             "@������������������������       �                     @                           Y@      �?             @������������������������       �                     �?������������������������       �                     @                           �S@"pc�
�?            �@@                           �N@���}<S�?             7@                           �L@r�q��?
             (@������������������������       �                     @                           @M@�q�q�?             @������������������������       �                     �?                            N@z�G�z�?             @������������������������       �                     @                          �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@!       $                    @M@���Q��?             $@"       #                    �K@���Q��?             @������������������������       �                      @������������������������       �                     @%       &                   �T@z�G�z�?             @������������������������       �                     �?������������������������       �                     @(       �                   @W@�HP��a�?�            pt@)       h                   @L@ z,m���?�             s@*       e                    �R@��<nd�?�            @k@+       d                    @O@Dw�&��?�            �j@,       C                    �J@|T(W�j�?f            �d@-       @                    @J@�? Da�?&            �O@.       ?                    �H@4և����?#             L@/       <                    @H@      �?             D@0       ;                    �G@�#-���?            �A@1       2                   �B@ȵHPS!�?             :@������������������������       �                     �?3       4                    �F@HP�s��?             9@������������������������       �        	             0@5       6                   �F@�<ݚ�?             "@������������������������       �                     @7       8                   @H@      �?             @������������������������       �                     �?9       :                    @G@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@=       >                    J@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@A       B                    E@և���X�?             @������������������������       �                     @������������������������       �                     @D       E                    @L@�:�]��?@            �Y@������������������������       �                    �A@F       W                    @M@t�U����?+            �P@G       H                    &@�+$�jP�?             ;@������������������������       �                     �?I       P                    �L@8�Z$���?             :@J       O                   �H@"pc�
�?             &@K       N                   @@@ףp=
�?             $@L       M                    :@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?Q       V                   @B@�r����?	             .@R       U                   �@@z�G�z�?             $@S       T                    =@      �?              @������������������������       �      �?             @������������������������       �                     @������������������������       �      �?              @������������������������       �                     @X       ]                    /@��(\���?             D@Y       Z                    '@      �?             @������������������������       �                      @[       \                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?^       _                    �M@�X�<ݺ?             B@������������������������       �                     *@`       a                   @E@���}<S�?             7@������������������������       �        	             &@b       c                   �F@r�q��?             (@������������������������       ��q�q�?             @������������������������       �                     "@������������������������       �                      I@f       g                    B@�q�q�?             @������������������������       �                     �?������������������������       �                      @i       �                   �R@
�GN��?>             V@j       k                    @F@���X�?(             L@������������������������       �                     "@l       �                   `R@(���@��?"            �G@m       n                   �L@���X�K�?             �F@������������������������       �                     �?o       p                   @M@���!pc�?             F@������������������������       �                     @q       t                     H@�z�G��?             D@r       s                   �Q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?u       �                    P@4�2%ޑ�?            �A@v       }                   @O@X�<ݚ�?             "@w       |                    �M@���Q��?             @x       {                   @N@      �?             @y       z                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?~       �                    �O@      �?             @       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @L@ȵHPS!�?             :@�       �                   `P@      �?              @������������������������       �                     �?�       �                    �K@����X�?             @�       �                    �H@r�q��?             @������������������������       �                      @�       �                     J@      �?             @������������������������       �      �?              @������������������������       �                      @������������������������       �                     �?�       �                     P@�X�<ݺ?
             2@������������������������       �                     $@�       �                    `P@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   `U@      �?             @@������������������������       �                     7@�       �                    V@�<ݚ�?             "@�       �                   �U@      �?             @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �I@�G��l��?             5@�       �                    �D@�q�q�?             .@�       �                    �B@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �X@�����H�?             "@������������������������       �                     @�       �                   `Y@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @L@0�����?�            pu@�       �                    �?��r�Z}�?�            �m@�       �                    @G@p��@���?0            @U@������������������������       �                     @@�       �                    �?���C��?             �J@������������������������       �                     <@�       �                    �G@�+e�X�?             9@������������������������       �                      @�       �                    A@�㙢�c�?             7@������������������������       �                     �?�       �                   `P@��2(&�?             6@������������������������       �                     (@�       �                    @I@�z�G��?             $@������������������������       �                     @������������������������       �                     @�       �                    @�=A�F�?]             c@�       �                   �J@~F�̫�?X            �a@�       �                    @G@�q�q�?             8@������������������������       �                     @�       �                    �G@�z�G��?             4@������������������������       �                     �?�       �                    @H@�����?             3@������������������������       �                     �?�       �                    �H@�E��ӭ�?
             2@������������������������       �                      @�       �                    �I@     ��?	             0@������������������������       �                     �?�       �                    �?������?             .@�       �                   �8@      �?              @������������������������       �                     @������������������������       �                     @�       �                   @H@؇���X�?             @�       �                    E@�q�q�?             @������������������������       �                     �?�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   @S@L�'�7��?I            @]@�       �                     B@z�G�z�?            �A@������������������������       �                      @�       �                    P@6YE�t�?            �@@������������������������       �                     2@�       �                    �?�q�q�?
             .@�       �                   `R@z�G�z�?             $@������������������������       �                      @�       �                    �E@      �?              @������������������������       �                     @�       �                    �H@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �G@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �\@������?2            �T@�       �                   �V@ ��WV�?0            �S@�       �                    V@�8��8��?             B@�       �                    @K@�IєX�?             A@�       �                    U@ 7���B�?             ;@������������������������       �                     0@�       �                    �B@�C��2(�?             &@�       �                    @@@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �T@؇���X�?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �      �?              @������������������������       �                     E@�       �                    �D@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �S@�eP*L��?             &@������������������������       �                     @�       �                    �B@      �?              @������������������������       �                     �?�       �                   �W@؇���X�?             @������������������������       �                     @�       �                   �Y@      �?             @������������������������       �                     �?������������������������       �                     @�       
      	             �?~|z����?F            �Z@�       	                   @��<b���?             7@�                         �D@�q�q�?
             .@                          �M@z�G�z�?             @������������������������       �                      @                        �7@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �?ףp=
�?             $@������������������������       �                     @                         �Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @      .                   @O@�!>�R�?8            �T@      #                   �M@t�F�}�?!            �I@                         �L@z�G�z�?             9@                         �?      �?              @������������������������       �                     @                        �U@�q�q�?             @������������������������       �                      @������������������������       �                     �?      "                  �V@������?             1@                         �?�	j*D�?             *@                         @M@�q�q�?             @                         H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?      !                   @z�G�z�?             $@                         @M@����X�?             @                        @P@      �?              @������������������������       �                     �?������������������������       �                     �?                          I@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @$      )                   @N@$��m��?             :@%      (                  �P@և���X�?             @&      '                  @K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @*      +                  @N@�����?	             3@������������������������       �                     (@,      -                   @؇���X�?             @������������������������       �                     @������������������������       �                     �?/      0                  @C@     ��?             @@������������������������       �                     @1      4                   �?�	j*D�?             :@2      3                  @J@r�q��?             @������������������������       �                     �?������������������������       �                     @5      B                  �T@��Q��?             4@6      A                   S@�E��ӭ�?             2@7      8                   �P@�q�q�?             .@������������������������       �                     @9      :                   �P@�q�q�?	             (@������������������������       �                     �?;      >                   @���|���?             &@<      =                  �K@և���X�?             @������������������������       �                     @������������������������       �                     @?      @                  �I@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @ri  trj  bh�h"h#K �rk  h%�rl  Rrm  (KMCKK�rn  hV�B0        t@     �y@     @Q@      t@      8@      D@      2@      *@      $@      (@              @      $@      @      @      �?              �?      @              @      @      �?      @      �?                      @      @               @      �?      @              @      �?              �?      @              @      ;@       @      5@       @      $@              @       @      @      �?              �?      @              @      �?      �?      �?                      �?              &@      @      @      @       @               @      @              �?      @      �?                      @     �F@     �q@     �A@     �p@      2@      i@      0@     �h@      0@     �b@       @     �K@      @     �I@      @     �A@      @      @@      @      7@      �?               @      7@              0@       @      @              @       @       @      �?              �?       @               @      �?                      "@       @      @              @       @                      0@      @      @      @                      @       @     �W@             �A@       @     �M@      @      6@      �?              @      6@       @      "@      �?      "@      �?      @              @      �?                      @      �?               @      *@       @       @      �?      @      �?      @              @      �?      �?              @      @     �B@      �?      @               @      �?      �?              �?      �?               @      A@              *@       @      5@              &@       @      $@       @      �?              "@              I@       @      �?              �?       @              1@     �Q@      .@     �D@              "@      .@      @@      *@      @@      �?              (@      @@              @      (@      <@      @      �?      @                      �?       @      ;@      @      @       @      @      �?      @      �?      �?              �?      �?                       @      �?              @      �?      �?      �?      �?                      �?       @              @      7@       @      @              �?       @      @      �?      @               @      �?      @      �?      �?               @      �?              �?      1@              $@      �?      @      �?                      @       @               @      >@              7@       @      @       @       @      �?      �?      �?                      �?      �?      �?              �?      �?                      @      $@      &@      $@      @       @      @       @                      @       @      �?      @              @      �?              �?      @                      @     `o@      W@      i@      B@     �S@      @      @@             �G@      @      <@              3@      @               @      3@      @              �?      3@      @      (@              @      @              @      @             �^@      >@      ]@      9@      $@      ,@      @              @      ,@              �?      @      *@      �?              @      *@               @      @      &@      �?              @      &@      @      @              @      @              �?      @      �?       @              �?      �?      �?      �?                      �?              @     �Z@      &@      <@      @               @      <@      @      2@              $@      @       @       @       @              @       @      @               @       @               @       @               @      @       @                      @     �S@      @     �R@      @     �@@      @      @@       @      :@      �?      0@              $@      �?      @      �?      @                      �?      @              @      �?      @      �?      @                      �?      @              �?      �?      E@              @      �?      @                      �?      @      @              @      @       @              �?      @      �?      @              @      �?              �?      @              I@      L@      2@      @      $@      @      �?      @               @      �?       @      �?                       @      "@      �?      @               @      �?       @                      �?       @              @@     �I@      ,@     �B@      @      4@      �?      @              @      �?       @               @      �?              @      *@      @      "@       @      �?      �?      �?              �?      �?              �?               @       @       @      @      �?      �?              �?      �?              �?      @      �?                      @              @              @      "@      1@      @      @      @      �?              �?      @                      @      @      *@              (@      @      �?      @                      �?      2@      ,@              @      2@       @      @      �?              �?      @              *@      @      *@      @      $@      @      @              @      @              �?      @      @      @      @      @                      @      @      �?              �?      @              @                       @ro  trp  bubhhubh)�rq  }rr  (hhh	h
hNhKhKhG        hh hNhJX��vhG        hNhG        h<Kh=Kh>h"h#K �rs  h%�rt  Rru  (KK�rv  hV�C              �?rw  trx  bhJhZhEC       ry  �rz  Rr{  h^Kh_h`Kh"h#K �r|  h%�r}  Rr~  (KK�r  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMAhkh"h#K �r�  h%�r�  Rr�  (KMA�r�  hr�B8F         :                    �?���
%�?�           ��@       /                   �U@Ҿ�q���?h             e@                           �?XΥf��?H            �^@                           8@��h!��?            �L@������������������������       �                      @                          @L@^(��I�?            �K@                            Q@؇���X�?             5@                           C@ףp=
�?
             4@	       
                   �A@����X�?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     *@������������������������       �                     �?                           @M@�!���?             A@                          �T@���Q��?	             .@                           �I@�eP*L��?             &@                          @R@z�G�z�?             @������������������������       �                      @                            E@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           R@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                           `P@�KM�]�?	             3@������������������������       �                     1@������������������������       �                      @       (                    @����?*            @P@                           A@XB���?$             M@������������������������       �                     �?        !                    �?0�)AU��?#            �L@������������������������       �                    �@@"       '                     I@ �q�q�?             8@#       $                    S@�����H�?             "@������������������������       �                     @%       &                    U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     .@)       *                    �M@����X�?             @������������������������       �                      @+       .                     P@���Q��?             @,       -                   �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @0       1                    �?`�q�0ܴ?             �G@������������������������       �                     ;@2       9                    @ףp=
�?             4@3       8                   @X@�����H�?             2@4       7                    �H@�<ݚ�?             "@5       6                     E@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                      @;       �                   �L@��\20�?i           ��@<       q                    �?�>���?�            �q@=       p                    �R@�8��8��?�            �i@>       O                    @L@���"F��?�            `i@?       @                    @I@X;��?8            @V@������������������������       �                     <@A       F                    �I@�.ߴ#�?'            �N@B       E                    E@���Q��?             @C       D                   �?@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @G       H                    @K@�h����?#             L@������������������������       �                     ?@I       N                    �K@`2U0*��?             9@J       K                    8@؇���X�?             @������������������������       �                     @L       M                   �F@      �?             @������������������������       �      �?              @������������������������       �                      @������������������������       �        
             2@P       ]                    @M@X�X\,��?M            �\@Q       V                    �L@8����?             7@R       U                   @@@      �?              @S       T                    :@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @W       X                    =@���Q��?
             .@������������������������       �                     @Y       \                   @B@"pc�
�?             &@Z       [                   �@@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     @^       g                   �E@���L��?<            �V@_       `                    �O@�h����?'             L@������������������������       �                     <@a       f                     P@h�����?             <@b       e                   �?@      �?              @c       d                    ;@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@h       o                   �G@؇���X�?            �A@i       j                   @F@�E��ӭ�?	             2@������������������������       �      �?             @k       l                    @O@d}h���?             ,@������������������������       �                      @m       n                     P@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     1@������������������������       �                     �?r       �                   �K@�J�j�?1            �S@s       t                    @G@�d�����?/             S@������������������������       �                     @u       ~                    �?@���?T�?,            �Q@v       }                     N@X�Cc�?             ,@w       x                   �:@X�<ݚ�?             "@������������������������       �                      @y       |                   �D@����X�?             @z       {                    �L@r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     �?������������������������       �                     @       �                    @�k�'7��?!            �L@�       �                     P@ZՏ�m|�?            �H@�       �                   �J@������?            �B@�       �                   �F@�FVQ&�?            �@@������������������������       �        	             1@�       �                    �M@      �?	             0@�       �                   �G@      �?              @������������������������       �                     �?�       �                    �J@؇���X�?             @�       �                   �I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �L@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �P@�q�q�?             (@������������������������       �                      @�       �                   �H@z�G�z�?             $@�       �                     R@�����H�?             "@������������������������       �                     @�       �                   �?@�q�q�?             @������������������������       �                     �?�       �                    F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �K@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    @L@d�w<h��?�            �q@�       �                    �?��s���?t            �g@�       �                    [@�iޤ��?*            �P@�       �                    @C@
��[��?)            @P@������������������������       �                     "@�       �                   `T@��X��?#             L@�       �                    T@�n_Y�K�?            �C@�       �                     E@�q�q�?             B@�       �                     D@���Q��?             @������������������������       ��q�q�?             @�       �                   �P@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @F@¦	^_�?             ?@������������������������       �                      @�       �                   �P@�û��|�?             7@�       �                   �O@ףp=
�?             $@������������������������       �                      @�       �                    �G@      �?              @������������������������       �                     �?������������������������       �                     @�       �                   �Q@�n_Y�K�?
             *@������������������������       �                     @�       �                   �R@X�<ݚ�?             "@�       �                   `R@���Q��?             @�       �                    @H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @K@      �?             @������������������������       �                      @�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �W@@�0�!��?
             1@������������������������       �                     (@�       �                   �X@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    @E@6�`��V�?J             _@������������������������       �                     A@�       �                    �?���Z�?3            �V@�       �                   �\@�r����?            �F@�       �                    @K@�Ra����?             F@�       �                   �S@`Jj��?             ?@�       �                   `R@r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �        
             3@�       �                    R@�θ�?             *@�       �                   �P@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �I@F�����?            �F@�       �                    @H@r�q��?             8@�       �                    @     ��?
             0@�       �                    �F@X�Cc�?             ,@������������������������       �                     @�       �                    Q@�eP*L��?             &@������������������������       �                      @�       �                   �R@X�<ݚ�?             "@������������������������       �                     @�       �                   @S@�q�q�?             @������������������������       �                      @�       �                    �G@      �?             @�       �                    T@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �S@      �?              @������������������������       �                     @�       �                    U@      �?             @������������������������       �                      @������������������������       �                      @�       �                    @��s����?             5@�       �                    @K@z�G�z�?             4@�       �                    �J@�<ݚ�?
             2@�       �                    @J@      �?              @�       �                    Y@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   `Q@�z�G��?             $@������������������������       �                     @�       �                   @S@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�                         �O@n�C���?>            �V@�       �                    �M@��
ц��?             *@������������������������       �                     @                          �?���Q��?             $@                        @M@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                        �R@�θ�?6            �S@                        �P@�S����?             C@                         �L@���N8�?             5@������������������������       �                     �?	                         �M@z�G�z�?             4@
                         @M@���Q��?             @������������������������       �                     @������������������������       �                      @                         �N@�r����?	             .@������������������������       �                     @                         �?      �?              @                        @P@؇���X�?             @                          P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                        `Q@�IєX�?             1@                         �?      �?              @������������������������       �                     @                         �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@      4                  �U@�z�G��?             D@      #                   �?�ՙ/�?             5@                         �S@z�G�z�?             @������������������������       �                      @!      "                  �T@�q�q�?             @������������������������       �                     �?������������������������       �                      @$      1                  `U@     ��?             0@%      ,                   �M@�q�q�?             (@&      +                   U@      �?             @'      (                   �?���Q��?             @������������������������       �                      @)      *                  �S@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?-      0                  �S@r�q��?             @.      /                   S@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @2      3                   �?      �?             @������������������������       �                     �?������������������������       �                     @5      8                   �L@���y4F�?             3@6      7                   Z@      �?             @������������������������       �                      @������������������������       �                      @9      @                   @�r����?
             .@:      ?                   Z@"pc�
�?             &@;      >                  �W@ףp=
�?             $@<      =                  `V@r�q��?             @������������������������       �                     @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMAKK�r�  hV�B       0s@     �z@     �^@     �G@     @S@     �F@      0@     �D@       @              ,@     �D@      @      2@       @      2@       @      @              @       @      �?              *@      �?              &@      7@      "@      @      @      @      �?      @               @      �?       @               @      �?              @       @      @                       @      @               @      1@              1@       @             �N@      @      L@       @              �?      L@      �?     �@@              7@      �?       @      �?      @              �?      �?              �?      �?              .@              @       @       @              @       @      �?       @      �?                       @       @             �F@       @      ;@              2@       @      0@       @      @       @      �?       @      �?                       @      @              "@               @              g@     �w@      D@     `n@      1@     `g@      0@     `g@      @     �U@              <@      @      M@       @      @       @      �?              �?       @                       @      �?     �K@              ?@      �?      8@      �?      @              @      �?      @      �?      �?               @              2@      *@     @Y@      @      0@      �?      @      �?      @              @      �?                      @      @      "@      @               @      "@       @      @              �?       @       @              @      @     @U@      �?     �K@              <@      �?      ;@      �?      @      �?       @               @      �?                      @              4@      @      >@      @      *@       @       @      @      &@               @      @      @      @                      @              1@      �?              7@      L@      4@      L@      @              .@      L@      @      "@      @      @               @      @       @      @      �?      @               @      �?              �?              @      $@     �G@       @     �D@      @     �@@       @      ?@              1@       @      ,@       @      @      �?              �?      @      �?       @      �?                       @              @               @       @       @       @                       @      @       @       @               @       @      �?       @              @      �?       @              �?      �?      �?      �?                      �?      �?               @      @       @                      @      @              b@      a@     @^@     �Q@      4@     �G@      2@     �G@              "@      2@      C@      .@      8@      (@      8@      @       @       @      �?      �?      �?              �?      �?              "@      6@               @      "@      ,@      �?      "@               @      �?      @      �?                      @       @      @      @              @      @      @       @      �?       @               @      �?               @              �?      @               @      �?      �?      �?                      �?      @              @      ,@              (@      @       @      @                       @       @             @Y@      7@      A@             �P@      7@     �C@      @     �C@      @      =@       @      $@       @      $@                       @      3@              $@      @      @      @      @                      @      @                      �?      <@      1@      &@      *@      "@      @      "@      @      @              @      @       @              @      @              @      @       @       @               @       @      �?       @               @      �?              �?                       @       @      @              @       @       @       @                       @      1@      @      0@      @      ,@      @      @      �?      @      �?      @                      �?      @              @      @      @               @      @              @       @               @              �?              8@     �P@      @      @              @      @      @      �?      @              @      �?              @              2@      N@      @      @@      @      0@      �?              @      0@       @      @              @       @               @      *@              @       @      @      �?      @      �?       @               @      �?                      @      �?              �?      0@      �?      @              @      �?      �?              �?      �?                      "@      (@      <@       @      *@      �?      @               @      �?       @      �?                       @      @      "@      @       @      @      @      @       @       @              �?       @               @      �?                      �?      �?      @      �?       @               @      �?                      @      @      �?              �?      @              @      .@       @       @       @                       @       @      *@       @      "@      �?      "@      �?      @              @      �?       @              @      �?                      @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ���EhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMwhkh"h#K �r�  h%�r�  Rr�  (KMw�r�  hr�BR         N       	             �?�r,��?�           ��@       C                   �U@�q����?h            �c@                          `P@��>4և�?L             \@                           �J@r�qG�?              H@                           �G@��2(&�?             6@������������������������       �                     @                          @C@     ��?             0@       	                   �A@���Q��?             @������������������������       �                     �?
                           �H@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     &@                           I@�n_Y�K�?             :@                           @      �?             4@                           �M@      �?
             0@������������������������       �                      @                           �?      �?              @                           �O@r�q��?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                          �A@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @       ,                    �K@     ��?,             P@       +                   �T@�q�q�?            �@@       $                    �?� �	��?             9@        #                    @H@�<ݚ�?             "@!       "                    �C@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @%       &                    �?      �?             0@������������������������       �                      @'       (                   �P@      �?              @������������������������       �                      @)       *                   �S@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @-       2                    S@f���M�?             ?@.       1                    Q@z�G�z�?             .@/       0                   �P@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     "@3       4                   �S@      �?             0@������������������������       �                     @5       B                    �O@�n_Y�K�?	             *@6       A                    @O@���!pc�?             &@7       <                    �N@�z�G��?             $@8       ;                   �U@����X�?             @9       :                    U@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @=       >                   `T@�q�q�?             @������������������������       �                     �??       @                    U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @D       K                    @O@dP-���?            �G@E       F                    @G@�(\����?             D@������������������������       �                     :@G       H                   �W@@4և���?             ,@������������������������       �                     &@I       J                   @X@�q�q�?             @������������������������       �                     �?������������������������       �                      @L       M                    X@և���X�?             @������������������������       �                     @������������������������       �                     @O       �                    �?�)	G!�?h           ��@P       �                    �M@B��h��?�            �u@Q       �                    @M@�q�q��?�             n@R       S                    @D@&��f���?�            `k@������������������������       �                     4@T       �                   @O@rLTAf�?y            �h@U       j                   @C@��ϻ�r�?P            ``@V       a                   �A@r�����?            �J@W       X                    @L@��(\���?             D@������������������������       �                     8@Y       `                    =@     ��?             0@Z       _                    :@      �?              @[       \                    5@r�q��?             @������������������������       �                     @]       ^                    8@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @b       c                    @G@��
ц��?             *@������������������������       �                     @d       g                   @B@      �?              @e       f                    @L@�q�q�?             @������������������������       �                      @������������������������       �                     �?h       i                    �J@z�G�z�?             @������������������������       �                     �?������������������������       �                     @k       t                   @I@$�q-�?3            �S@l       m                   �F@�(\����?             D@������������������������       �                     ,@n       s                   @G@ ��WV�?             :@o       r                    �H@�8��8��?
             (@p       q                    @F@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@u       v                    �E@�?�'�@�?             C@������������������������       �                     @w       �                    �H@     ��?             @@x       }                   �J@�q�q�?             "@y       z                    �F@�q�q�?             @������������������������       �                     �?{       |                    @G@      �?              @������������������������       �                     �?������������������������       �                     �?~       �                   �L@r�q��?             @       �                    @H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �M@���}<S�?             7@�       �                   �J@P���Q�?             4@�       �                    �K@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     &@�       �                   @N@�q�q�?             @�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �L@�l�]�N�?)             Q@�       �                   @Z@     ��?'             P@�       �                   �R@f�<�>��?$            �M@�       �                   `R@      �?             B@�       �                   �P@��}*_��?             ;@�       �                    P@�G�z��?             4@������������������������       �                     �?�       �                   �P@D�n�3�?             3@�       �                    @K@b�2�tk�?
             2@�       �                    �I@8�Z$���?             *@�       �                   `P@�q�q�?             @������������������������       �                     �?�       �                    @F@���Q��?             @������������������������       �                      @�       �                    �G@�q�q�?             @������������������������       �                     �?�       �                    �H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   `Q@؇���X�?             @�       �                    @I@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �K@�����H�?             "@������������������������       �                     @������������������������       �z�G�z�?             @�       �                   �W@��+7��?             7@�       �                    �J@8�Z$���?	             *@������������������������       �                     "@�       �                   �R@      �?             @������������������������       �                     �?�       �                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �X@���Q��?             $@�       �                    X@�q�q�?             @�       �                    �G@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    K@�G��l��?             5@������������������������       �                     @�       �                   �M@      �?             0@������������������������       �                      @�       �                   �O@և���X�?             ,@������������������������       �                      @�       �                   �P@�q�q�?             (@������������������������       �z�G�z�?             @�       �                   `S@և���X�?             @������������������������       �                      @�       �                   �U@z�G�z�?             @������������������������       �                     @�       �                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    `P@�:�H:�?E            @[@�       �                   @E@�o��gn�?2            �T@�       �                    @O@г�wY;�?             A@�       �                    �N@�8��8��?             (@������������������������       �                     @�       �                    3@r�q��?             @�       �                    $@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@�       �                   @G@�����?            �H@�       �                    @O@�n_Y�K�?             *@�       �                   �F@      �?              @������������������������       �      �?             @������������������������       �                     @�       �                     P@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   @M@4?,R��?             B@�       �                    �O@P���Q�?             4@������������������������       �                     *@�       �                     P@؇���X�?             @�       �                   �K@      �?             @�       �                   �I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                     P@      �?             0@�       �                   �N@�C��2(�?
             &@������������������������       �                     �?������������������������       �        	             $@�       �                   �R@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     :@�       >                   �L@��\20�?�            @l@�                          N@ ]�к��?b             b@�       �                    �G@8�A�0��?             6@������������������������       �                     @�       �                   �D@�\��N��?             3@�       �                    �J@�q�q�?             (@�       �                    @I@�����H�?             "@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   @H@����X�?             @������������������������       �                     @�                         �J@�q�q�?             @                          �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?      /                  �U@,���i�?S            �^@      &                   T@$gv&��?*            �M@                         �E@ZՏ�m|�?#            �H@������������������������       �        
             1@      %                   @      �?             @@	                         �I@��a�n`�?             ?@
                         �G@���Q��?	             $@                         @F@�q�q�?             @                         R@      �?              @������������������������       �                     �?������������������������       �                     �?                        �R@      �?             @                         �F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         �?      �?             @������������������������       �                     �?                        �S@�q�q�?             @������������������������       �                      @������������������������       �                     �?                         �?؇���X�?             5@                         Q@$�q-�?
             *@������������������������       �                      @                         R@z�G�z�?             @������������������������       �                     �?������������������������       �                     @      $                  @S@      �?              @       #                   �K@      �?             @!      "                  `Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?'      .                   @���Q��?             $@(      )                   �B@      �?              @������������������������       �                     �?*      +                   @K@؇���X�?             @������������������������       �                     @,      -                  �T@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @0      1                   �G@     �?)             P@������������������������       �                     E@2      7                   �I@��2(&�?             6@3      4                   �?���Q��?             @������������������������       �                     �?5      6                  �W@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?8      =                   @K@�IєX�?
             1@9      <                   �?r�q��?             @:      ;                   �J@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@?      L                   �?(Q��h�?1            @T@@      E                   �N@�X����?             6@A      D                  @T@�eP*L��?             &@B      C                  @H@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @F      I                    Q@"pc�
�?             &@G      H                  �K@      �?              @������������������������       �                     @������������������������       �                     �?J      K                  �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?M      j                   �P@�ݜ����?%            �M@N      e                   @v ��?            �E@O      d                   @P@�xGZ���?            �A@P      Y                  �L@�'�=z��?            �@@Q      T                   @@�q�q�?             2@R      S                   @M@z�G�z�?             @������������������������       �                     �?������������������������       �                     @U      X                   �M@8�Z$���?             *@V      W                   H@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @Z      c                    O@������?             .@[      b                  �W@d}h���?             ,@\      a                  @R@8�Z$���?             *@]      ^                  �O@����X�?             @������������������������       �                     @_      `                   �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @f      g                  �L@      �?              @������������������������       �                     @h      i                   U@z�G�z�?             @������������������������       �                     @������������������������       �                     �?k      v                   S@     ��?             0@l      u                   P@d}h���?
             ,@m      n                    Q@�q�q�?             "@������������������������       �                     @o      p                   D@      �?             @������������������������       �                      @q      t                   @      �?             @r      s                   �R@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMwKK�r�  hV�Bp       �t@     Py@     �[@      H@      Q@      F@     �A@      *@      3@      @      @              *@      @       @      @              �?       @       @      �?              �?       @      &@              0@      $@      $@      $@      @      $@               @      @       @      @      �?      @               @      �?              �?       @              �?      �?      �?                      �?      @              @             �@@      ?@      6@      &@      ,@      &@       @      @       @      @              @       @                      @      (@      @       @              @      @               @      @       @      @                       @       @              &@      4@      @      (@      @      @              @      @                      "@       @       @      @              @       @      @       @      @      @       @      @       @       @               @       @                      @      �?       @              �?      �?      �?      �?                      �?              �?       @             �E@      @     �C@      �?      :@              *@      �?      &@               @      �?              �?       @              @      @              @      @             @k@     Pv@     �P@     �q@     �K@      g@     �F@     �e@              4@     �F@     @c@      0@     �\@      $@     �E@      @     �B@              8@      @      *@      @      @      �?      @              @      �?       @      �?                       @       @                       @      @      @      @               @      @      �?       @               @      �?              �?      @      �?                      @      @      R@      �?     �C@              ,@      �?      9@      �?      &@      �?      @              @      �?                       @              ,@      @     �@@              @      @      ;@      @      @       @      �?      �?              �?      �?              �?      �?              �?      @      �?       @               @      �?                      @       @      5@      �?      3@      �?       @               @      �?                      &@      �?       @      �?      �?              �?      �?                      �?      =@     �C@      =@     �A@      8@     �A@      2@      2@      $@      1@      "@      &@      �?               @      &@      @      &@       @      &@       @      @              �?       @      @               @       @      �?      �?              �?      �?              �?      �?                      @      @              �?              �?      @      �?      @      �?                      @              @       @      �?      @              @      �?      @      1@       @      &@              "@       @       @              �?       @      �?       @                      �?      @      @      @       @       @       @       @                       @       @                      @      @                      @      $@      &@              @      $@      @       @               @      @               @       @      @      @      �?      @      @               @      @      �?      @              �?      �?              �?      �?              &@     �X@      &@      R@      �?     �@@      �?      &@              @      �?      @      �?       @               @      �?                      @              6@      $@     �C@      @       @       @      @       @       @              @      @       @      @                       @      @      ?@      �?      3@              *@      �?      @      �?      @      �?      �?              �?      �?                       @              @      @      (@      �?      $@      �?                      $@      @       @      @                       @              :@      c@     �R@     @]@      <@      "@      *@              @      "@      $@      @       @      �?       @      �?      @      �?                      @              @      @              @       @      @              �?       @      �?      �?      �?                      �?              �?      [@      .@     �G@      (@     �D@       @      1@              8@       @      8@      @      @      @      @       @      �?      �?      �?                      �?      @      �?      �?      �?      �?                      �?       @               @       @      �?              �?       @               @      �?              2@      @      (@      �?       @              @      �?              �?      @              @       @       @       @       @      �?       @                      �?              �?      @                      �?      @      @      @       @              �?      @      �?      @               @      �?              �?       @                       @     �N@      @      E@              3@      @      @       @              �?      @      �?       @      �?      �?              0@      �?      @      �?      @      �?      @                      �?      �?              &@             �A@      G@      @      .@      @      @      @      �?              �?      @                      @       @      "@      �?      @              @      �?              �?       @               @      �?              <@      ?@      7@      4@      3@      0@      1@      0@      @      (@      @      �?              �?      @               @      &@       @      @       @                      @              @      &@      @      &@      @      &@       @      @       @      @              �?       @               @      �?              @                      �?              �?       @              @      @              @      @      �?      @                      �?      @      &@      @      &@      @      @              @      @      @               @      @      �?       @      �?       @                      �?      �?                      @       @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ:9)bhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMhkh"h#K �r�  h%�r�  Rr�  (KM�r�  hr�BX>         :                    �?T8���?�           ��@       -                   �T@�<ݚ��?_             b@                           @H@�
�G�?9             V@                           �?�C��2(�?             6@                           �D@      �?              @������������������������       �                     �?                           �G@؇���X�?             @������������������������       �                     @	       
                   �A@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@       "                    �?8�A�0��?+            �P@                           �J@և���X�?            �A@                           �I@����X�?             ,@                           @I@      �?              @������������������������       �      �?             @                          �F@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       !                    �P@���N8�?             5@                           @L@�S����?             3@������������������������       �                     @                          �N@d}h���?             ,@                           �O@      �?             @������������������������       �                      @������������������������       �                      @                           �O@ףp=
�?             $@������������������������       �                     @                           @R@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @#       $                    C@��a�n`�?             ?@������������������������       �                      @%       &                    �?д>��C�?             =@������������������������       �        
             .@'       (                   @O@X�Cc�?	             ,@������������������������       �                     @)       *                   @R@      �?              @������������������������       �                     @+       ,                    T@      �?             @������������������������       �                     @������������������������       �                     �?.       9                   �W@h�����?&             L@/       0                    �N@�FVQ&�?            �@@������������������������       �                     7@1       8                    @P@z�G�z�?             $@2       7                    @O@����X�?             @3       4                    U@r�q��?             @������������������������       �                     @5       6                   �U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     7@;       �                    �?2� J��?p           p�@<       �                    P@h~��M�?�            �t@=       n                   @C@X	
bi��?�            @n@>       ?                    �D@ܔQ|ӭ�?H            �[@������������������������       �                     �?@       m                    �R@�~i��?G            @[@A       D                    �I@d/
k�?F             [@B       C                     I@      �?             (@������������������������       �                     "@������������������������       �                     @E       d                    @O@�8��8��??             X@F       G                    @K@     ��?+             P@������������������������       �                     "@H       Q                    .@X�;�^o�?$            �K@I       J                    �L@���!pc�?             &@������������������������       �                     @K       L                    �M@      �?              @������������������������       �                     �?M       N                    '@����X�?             @������������������������       �                     @O       P                    �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @R       Y                   �A@�C��2(�?             F@S       T                    �L@      �?             @@������������������������       �                     (@U       X                    @M@P���Q�?             4@V       W                    =@      �?              @������������������������       �      �?              @������������������������       �                     @������������������������       �                     (@Z       ]                     L@      �?
             (@[       \                   @B@      �?             @������������������������       ��q�q�?             @������������������������       �                     �?^       c                    �M@      �?              @_       `                    �L@z�G�z�?             @������������������������       �                      @a       b                   @B@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @e       f                   �>@      �?             @@������������������������       �        
             2@g       l                     P@@4և���?
             ,@h       i                    �O@r�q��?             @������������������������       �                     @j       k                   �?@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?o       p                    @H@���7�?T            �`@������������������������       �                    �B@q       x                   �K@8v�YeK�??            �W@r       s                    �O@�"w����?2             S@������������������������       �        )             N@t       u                   �J@      �?	             0@������������������������       �                     ,@v       w                   @K@      �?              @������������������������       �                     �?������������������������       �                     �?y       z                    �I@�d�����?             3@������������������������       �                     @{       |                   @L@      �?             0@������������������������       �                     @}       �                    N@r�q��?             (@~                           @M@�<ݚ�?             "@������������������������       �                     @�       �                   �L@���Q��?             @������������������������       �                     �?�       �                   @M@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   @W@�^�����?>            �U@�       �                    @D@      �?.             P@������������������������       �                     (@�       �                   �R@�	j*D�?'             J@�       �                    @H@     ��?             @@�       �                    �F@      �?              @�       �                   �Q@      �?             @������������������������       �                      @�       �                   `R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    R@      �?             8@�       �                    �O@��s����?             5@�       �                   �P@�S����?             3@�       �                   �P@���!pc�?
             &@�       �                    �K@z�G�z�?	             $@������������������������       �                     @�       �                    �L@���Q��?             @������������������������       �                     �?�       �                    @M@      �?             @������������������������       �                     �?�       �                    �M@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `R@�q�q�?             @������������������������       �                     �?�       �                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    T@R���Q�?             4@������������������������       �                     (@�       �                   `T@      �?              @������������������������       �                      @�       �                   `U@r�q��?             @������������������������       �                     @�       �                   �U@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �W@�eP*L��?             6@������������������������       �                     @�       �                    �D@p�ݯ��?             3@������������������������       �                     @�       �                   �Y@      �?
             ,@�       �                    Y@���Q��?             $@�       �                    X@      �?              @�       �                    �G@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                     K@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �K@�E�-���?�            `p@�       �                    �?�z�G��?&            �Q@�       �                   �8@�G�z��?             4@������������������������       �                     @�       �                     N@������?             .@�       �                   �F@�8��8��?             (@������������������������       �                      @�       �                    �K@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @z�G�z�?             I@�       �                   �1@�GN�z�?             F@�       �                    �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @I@� ��1�?            �D@�       �                   �D@�S����?             C@�       �                   �;@�C��2(�?
             6@�       �                     N@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     .@�       �                    �K@      �?	             0@������������������������       �                      @�       �                    F@؇���X�?             ,@������������������������       �                     �?�       �                     P@$�q-�?             *@������������������������       �                     "@�       �                    �Q@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�                          @r�q�?p             h@�       �                    S@b�h�d.�?f            �e@�       �                    P@����>�?(            �R@������������������������       �                     9@�       �                    �?ڡR����?            �H@�       �                    �B@      �?             8@������������������������       �                      @�       �                    @K@"pc�
�?             6@������������������������       �                     &@�       �                    �L@���|���?             &@�       �                     L@և���X�?             @������������������������       �                     �?�       �                   �P@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �F@� �	��?             9@������������������������       �                     @�       �                   �R@�<ݚ�?	             2@�       �                   �P@ףp=
�?             $@�       �                   `P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @H@      �?              @������������������������       �                     @������������������������       �                     @                          �?ܴD��?>            @Y@                        `\@ �#�Ѵ�?            �E@������������������������       �                     D@                         �D@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �H@\-��p�?#             M@������������������������       �                     9@                         �P@r٣����?            �@@	                         �O@������?             >@
                         Y@>���Rp�?             =@                        �T@8�Z$���?             :@                         T@����X�?             @������������������������       �                     @������������������������       �                      @                        �U@�KM�]�?             3@������������������������       �                      @                         �L@"pc�
�?             &@                        �V@ףp=
�?             $@������������������������       �      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @                         �N@ҳ�wY;�?
             1@                         X@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hV�B�       �t@     @y@     @\@      ?@     �M@      =@      4@       @      @       @              �?      @      �?      @              �?      �?              �?      �?              ,@             �C@      ;@      .@      4@      $@      @      @      @      @      �?      �?      @      �?                      @      @              @      0@      @      0@              @      @      &@       @       @       @                       @      �?      "@              @      �?      @              @      �?               @              8@      @               @      8@      @      .@              "@      @      @              @      @              @      @      �?      @                      �?      K@       @      ?@       @      7@               @       @      @       @      @      �?      @              �?      �?              �?      �?                      �?      @              7@              k@     Pw@     �F@     �q@      3@     �k@      *@     @X@      �?              (@     @X@      &@     @X@      @      "@              "@      @               @      V@      @     �L@              "@      @      H@      @       @              @      @      @      �?               @      @              @       @      �?              �?       @              @      D@      �?      ?@              (@      �?      3@      �?      @      �?      �?              @              (@      @      "@       @       @       @      �?              �?      �?      @      �?      @               @      �?       @      �?      �?              �?              @      �?      ?@              2@      �?      *@      �?      @              @      �?      �?      �?                      �?               @      �?              @     �_@             �B@      @     @V@      �?     �R@              N@      �?      .@              ,@      �?      �?      �?                      �?      @      ,@      @               @      ,@              @       @      $@       @      @              @       @      @      �?              �?      @              @      �?                      @      :@      N@      0@      H@              (@      0@      B@      *@      3@      @      �?      @      �?       @              �?      �?              �?      �?              @              @      2@      @      1@      @      0@      @       @       @       @              @       @      @      �?              �?      @              �?      �?       @      �?      �?              �?      �?                       @      �?      �?      �?                      �?       @      �?      �?              �?      �?      �?                      �?      @      1@              (@      @      @       @              �?      @              @      �?       @      �?                       @      $@      (@      @              @      (@              @      @      @      @      @      @      @       @      @       @                      @       @                       @      @      �?      @                      �?     �e@     �V@      5@     �H@      &@      "@              @      &@      @      &@      �?       @              @      �?      @                      �?              @      $@      D@      $@      A@       @      �?              �?       @               @     �@@      @      @@       @      4@       @      @       @                      @              .@      @      (@       @               @      (@      �?              �?      (@              "@      �?      @      �?                      @       @      �?              �?       @                      @     �b@     �D@      b@      >@      K@      4@      9@              =@      4@      2@      @               @      2@      @      &@              @      @      @      @              �?      @      @      @                      @      @              &@      ,@      @              @      ,@      �?      "@      �?      �?              �?      �?                       @      @      @      @                      @     �V@      $@     �D@       @      D@              �?       @      �?                       @      I@       @      9@              9@       @      6@       @      6@      @      6@      @      @       @      @                       @      1@       @       @              "@       @      "@      �?      @      �?      @                      �?              @              �?      @              @      &@      �?      &@              &@      �?              @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�BHzhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjMihkh"h#K �r�  h%�r�  Rr�  (KMi�r�  hr�B�N         <                    �?�[��N�?�           ��@       %                    �?V������?]            �b@                          �T@�w��#��?%             I@                           `P@��Q���?             D@                           �J@�I�w�"�?             C@                           Q@      �?             0@                          �P@z�G�z�?             $@                          �N@����X�?             @	       
                    �H@r�q��?             @������������������������       �                     @                           @I@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          @R@�q�q�?             @������������������������       �                     @������������������������       �                      @                            N@��2(&�?             6@������������������������       �                     *@                           S@�q�q�?             "@                          �G@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @       $                   �V@���Q��?	             $@                           @M@      �?              @������������������������       �                     @                           �N@      �?             @������������������������       �                     �?        !                    U@�q�q�?             @������������������������       �                     �?"       #                   �U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @&       1                    �J@�+�$f��?8            �X@'       (                    �?XB���?!             M@������������������������       �                     >@)       *                   �S@@4և���?             <@������������������������       �        	             4@+       ,                    @G@      �?              @������������������������       �                     @-       .                   �T@���Q��?             @������������������������       �                     �?/       0                   �V@      �?             @������������������������       �                     @������������������������       �                     �?2       ;                    @R���Q�?             D@3       4                   �C@      �?             B@������������������������       �                     @5       6                    �? 	��p�?             =@������������������������       �                     $@7       :                   �J@�KM�]�?
             3@8       9                    �R@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     .@������������������������       �                     @=       �                   @L@�ΫY�^�?j           P�@>       K                    �D@�����U�?�            0r@?       D                   @C@      �?             0@@       C                    �?�<ݚ�?             "@A       B                    �C@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @E       F                    �B@؇���X�?             @������������������������       �                     @G       H                    H@�q�q�?             @������������������������       �                     �?I       J                    �C@      �?              @������������������������       �                     �?������������������������       �                     �?L       �                   �I@�h�>(�?�            0q@M       n                    @K@�*/�8V�?�            `m@N       c                    @J@��a�2��?-             R@O       P                   �:@�r����?            �F@������������������������       �                     (@Q       b                    �I@"pc�
�?            �@@R       [                    �H@d}h���?             <@S       T                   �;@��2(&�?             6@������������������������       �                     �?U       V                    �?�����?             5@������������������������       �        
             *@W       X                   �C@      �?              @������������������������       �                     @Y       Z                    @G@�q�q�?             @������������������������       �                      @������������������������       �                     �?\       a                    �?      �?             @]       ^                    @I@      �?             @������������������������       �                     �?_       `                    E@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @d       i                    �?������?             ;@e       h                    �J@�����?             5@f       g                   �A@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             2@j       k                    �?r�q��?             @������������������������       �                      @l       m                   @F@      �?             @������������������������       �                     �?������������������������       �                     @o       �                    �Q@�u�w�u�?e            `d@p       �                    �?Х-��ٹ?\            �b@q       t                    @H��ԛ�?I            �]@r       s                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?u       v                    6@XB���?G             ]@������������������������       �                     8@w       z                   �7@�nkK�?;             W@x       y                     L@      �?              @������������������������       �                     �?������������������������       �                     �?{       �                    �K@(;L]n�?9            �V@|       }                   �?@      �?             @������������������������       �                     �?~                          @B@�q�q�?             @������������������������       �      �?              @������������������������       �                     �?�       �                   �A@ qP��B�?5            �U@������������������������       �                     >@�       �                   @B@h�����?$             L@�       �                    �M@      �?              @������������������������       �                     �?������������������������       �                     @�       �                   �F@@��8��?              H@������������������������       �                     <@�       �                   @G@P���Q�?             4@�       �                     P@ףp=
�?             $@�       �                    @O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �                    <@��a�n`�?             ?@�       �                    :@�q�q�?             "@�       �                   �0@z�G�z�?             @�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     6@�       �                   �C@�	j*D�?	             *@������������������������       �                     @�       �                    �?      �?              @������������������������       �                      @�       �                    �R@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �K@��Q��?             D@�       �                   @J@8�Z$���?             *@������������������������       �                     @�       �                   �J@      �?              @�       �                    @G@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �I@r�q��?             @�       �                    �G@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   @J@X�<ݚ�?             ;@�       �                    @L@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   @K@�<ݚ�?
             2@�       �                    �L@X�<ݚ�?             "@������������������������       �                     @�       �                    �?r�q��?             @�       �                   �J@�q�q�?             @������������������������       �                     �?�       �                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       0                   @L@���Zհ�?�            pr@�                         `U@���ٕ�?|            `h@�                           �K@)b���?B            �Z@�       �                    �?b*0t��?A            �Y@�       �                    @I@��h!��?!            �L@�       �                    Q@<���D�?            �@@�       �                    �E@������?
             .@������������������������       �                     @�       �                   `P@���|���?             &@������������������������       �                     @�       �                    �G@      �?              @������������������������       �                     @�       �                    �H@z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �        
             2@�       �                   �R@      �?             8@�       �                   �Q@D�n�3�?
             3@�       �                   @P@�n_Y�K�?             *@�       �                    O@�q�q�?             @�       �                   �M@�q�q�?             @������������������������       �                     �?�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �P@؇���X�?             @�       �                    @K@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �S@z�G�z�?             @�       �                    @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @K@�I� �?              G@�       �                    R@��Q���?             D@�       �                    �B@��2(&�?             6@������������������������       �                      @�       �                    @G@P���Q�?             4@�       �                    @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     $@�       �                   `T@X�<ݚ�?             2@�       �                    T@      �?             0@�       �                    @G@�q�q�?	             (@�       �                   �R@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                     J@z�G�z�?             @������������������������       �                     @�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @E@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    R@�q�q�?             @�       �                   �N@z�G�z�?             @�       �                   @M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @      /                   @K@�7�A�?:             V@                         �F@������?6            @T@                         �?j�q����?              I@                        �X@      �?	             (@                        @V@���Q��?             $@������������������������       �                     �?      	                   W@X�<ݚ�?             "@������������������������       �                     �?
                        �W@      �?              @������������������������       �                      @                         �D@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @                        `Z@�˹�m��?             C@                        �U@XB���?             =@                         �C@z�G�z�?             @                         @@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     8@                         @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @      (                   �I@���@M^�?             ?@      #                   X@     ��?             0@                         �?�q�q�?             "@������������������������       �                     @      "                   W@���Q��?             @       !                    H@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @������������������������       �                     �?$      %                   �G@և���X�?             @������������������������       �                      @&      '                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @)      .                  @[@z�G�z�?
             .@*      -                   �?$�q-�?	             *@+      ,                  �U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                      @������������������������       �                     @1      <                  �O@� �	��?;             Y@2      7                  @M@$��m��?             :@3      6                  �L@��
ц��?             *@4      5                    M@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @8      ;                   �?8�Z$���?             *@9      :                   N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@=      L                   S@�r*e���?-            �R@>      E                   �?��<b���?             G@?      D                   �M@ףp=
�?             >@@      C                  �P@�q�q�?             "@A      B                   @M@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     @������������������������       �                     5@F      G                  �Q@     ��?             0@������������������������       �                     @H      K                   �M@ףp=
�?             $@I      J                   �L@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @M      V                   �?��>4և�?             <@N      Q                  �W@      �?              @O      P                   �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?R      S                   @M@z�G�z�?             @������������������������       �                     @T      U                   �M@      �?              @������������������������       �                     �?������������������������       �                     �?W      X                   �L@�z�G��?             4@������������������������       �                     @Y      h                  �W@ҳ�wY;�?             1@Z      ]                   @M@d}h���?	             ,@[      \                  �T@      �?              @������������������������       �                     �?������������������������       �                     �?^      g                   �P@r�q��?             (@_      d                   �O@"pc�
�?             &@`      a                  �U@؇���X�?             @������������������������       �                     @b      c                  @V@      �?             @������������������������       �                     �?������������������������       �                     @e      f                  �T@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMiKK�r�  hV�B�       �s@     Pz@      Z@      F@      1@     �@@      &@      =@      "@      =@      @      $@       @       @       @      @      �?      @              @      �?       @      �?      �?              �?      �?                      @      @       @      @                       @      @      3@              *@      @      @      �?      @      �?                      @       @               @              @      @      @       @      @               @       @              �?       @      �?      �?              �?      �?              �?      �?                       @     �U@      &@      L@       @      >@              :@       @      4@              @       @      @              @       @              �?      @      �?      @                      �?      ?@      "@      ;@      "@              @      ;@       @      $@              1@       @       @       @               @       @              .@              @              j@     �w@     �G@     �n@       @       @      @       @       @       @               @       @              @              �?      @              @      �?       @              �?      �?      �?      �?                      �?     �C@     �m@      9@     @j@      *@     �M@      @     �C@              (@      @      ;@      @      6@      @      3@      �?               @      3@              *@       @      @              @       @      �?       @                      �?      @      @      �?      @              �?      �?       @      �?                       @       @                      @      @      4@       @      3@       @      �?              �?       @                      2@      @      �?       @              @      �?              �?      @              (@     �b@       @     �a@      @     �\@      �?       @               @      �?              @      \@              8@      @      V@      �?      �?              �?      �?              @     �U@      �?      @              �?      �?       @      �?      �?              �?       @      U@              >@       @      K@      �?      @      �?                      @      �?     �G@              <@      �?      3@      �?      "@      �?      @              @      �?                      @              $@      @      <@      @      @      �?      @      �?      �?              �?      �?                      @       @       @       @                       @              6@      @      "@              @      @      @               @      @       @      @                       @      ,@      :@       @      &@              @       @      @      �?      �?      �?                      �?      �?      @      �?       @               @      �?                      @      (@      .@       @      �?              �?       @              @      ,@      @      @      @              �?      @      �?       @              �?      �?      �?              �?      �?                      @              "@     @d@     �`@     �]@     @S@     �I@      L@     �G@      L@      0@     �D@      @      =@      @      &@              @      @      @              @      @      @      @              �?      @               @      �?       @              2@      (@      (@      &@       @      @       @      @       @      �?       @              �?      �?      �?              �?      �?              @              �?      @      �?      @              @      �?                      �?      @              �?      @      �?       @               @      �?                       @      ?@      .@      =@      &@      3@      @               @      3@      �?      "@      �?      "@                      �?      $@              $@       @       @       @      @      @      @      �?              �?      @              �?      @              @      �?      �?      �?                      �?      �?      @      �?                      @       @               @      @      �?      @      �?      �?              �?      �?                      @      �?              @             �P@      5@      N@      5@     �D@      "@      @      @      @      @      �?              @      @              �?      @      @       @              @      @              @      @                       @     �A@      @      <@      �?      @      �?      �?      �?      �?                      �?      @              8@              @       @      @                       @      3@      (@      @      "@      @      @              @      @       @      @      �?      �?               @      �?              �?      @      @               @      @      �?              �?      @              (@      @      (@      �?      �?      �?      �?                      �?      &@                       @      @              F@      L@      1@      "@      @      @      @      �?              �?      @                      @      &@       @      �?       @      �?                       @      $@              ;@     �G@      $@      B@      @      ;@      @      @      @       @              �?      @      �?              @              5@      @      "@      @              �?      "@      �?      @              @      �?                      @      1@      &@      @      @       @      �?       @                      �?      �?      @              @      �?      �?      �?                      �?      ,@      @      @              &@      @      &@      @      �?      �?      �?                      �?      $@       @      "@       @      @      �?      @              @      �?              �?      @              @      �?      @                      �?      �?                      @r�  tr�  bubhhubehhub.